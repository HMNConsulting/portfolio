<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<!-- Created with Inkscape (http://www.inkscape.org/) -->

<svg
   version="1.1"
   id="svg2340"
   width="1056"
   height="1632"
   viewBox="0 0 1056 1632"
   sodipodi:docname="header-bg.sv"
   inkscape:version="1.2.2 (732a01da63, 2022-12-09)"
   xmlns:inkscape="http://www.inkscape.org/namespaces/inkscape"
   xmlns:sodipodi="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd"
   xmlns:xlink="http://www.w3.org/1999/xlink"
   xmlns="http://www.w3.org/2000/svg"
   xmlns:svg="http://www.w3.org/2000/svg">
  <defs
     id="defs2344">
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath2354">
      <path
         d="m 455,1787 4,4 h 8169 l -2975,-4 h 2979 l -4,4 v 1925 l 12,-1929 v 1917 l 3558,12 H 8628 l 12,-12 h 3563 v 7 l -5,5 v 15212 l 5,-6343 v 6348 l -5,-5 H 459 l 4896,5 H 454 l 5,-5 V 1791 l -5,7145 V 1787 h 1"
         id="path2352" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath4082">
      <path
         d="m 455,1787 4,4 h 8169 l -2975,-4 h 2979 l -4,4 v 1925 l 12,-1929 v 1917 l 3558,12 H 8628 l 12,-12 h 3563 v 7 l -5,5 v 15212 l 5,-6343 v 6348 l -5,-5 H 459 l 4896,5 H 454 l 5,-5 V 1791 l -5,7145 V 1787 h 1"
         id="path4080" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath4090">
      <path
         d="m 455,1787 4,4 h 8169 l -2975,-4 h 2979 l -4,4 v 1925 l 12,-1929 v 1917 l 3558,12 H 8628 l 12,-12 h 3563 v 7 l -5,5 v 15212 l 5,-6343 v 6348 l -5,-5 H 459 l 4896,5 H 454 l 5,-5 V 1791 l -5,7145 V 1787 h 1"
         id="path4088" />
    </clipPath>
    <mask
       maskUnits="userSpaceOnUse"
       x="0"
       y="0"
       width="1"
       height="1"
       id="mask4094">
      <image
         width="1"
         height="1"
         style="image-rendering:optimizeSpeed"
         preserveAspectRatio="none"
         xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAADMAAAAzCAAAAAAfym/2AAAAAXNCSVQI5gpbmQAAALZJREFUSIntls0OhCAQg1ve/53Zg0aGrfx0TMwelgMy2o8yxMAQ2moXUb7LmyoS0XzFN4SqYjQARBfGM6RTttECCdKyjbRW1hKZlZYLQ7+9MALW2q7Ji2XTzCyEQLFd7HyAmmAyPqhJH3sLwAzjIy/t25/5dSbzvyV8mMtH77E1k/FxG33mOBPthAhYJylx5mM6mfkwWCTuuU2I3WMH0rve2IdndcicGtQ7E2pcV42wRf2m1I3gA/WBHU9CSSKCAAAAAElFTkSuQmCC"
         id="image4096" />
    </mask>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath4112">
      <path
         d="m 455,1787 4,4 h 8169 l -2975,-4 h 2979 l -4,4 v 1925 l 12,-1929 v 1917 l 3558,12 H 8628 l 12,-12 h 3563 v 7 l -5,5 v 15212 l 5,-6343 v 6348 l -5,-5 H 459 l 4896,5 H 454 l 5,-5 V 1791 l -5,7145 V 1787 h 1"
         id="path4110" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath4120">
      <path
         d="m 455,1787 4,4 h 8169 l -2975,-4 h 2979 l -4,4 v 1925 l 12,-1929 v 1917 l 3558,12 H 8628 l 12,-12 h 3563 v 7 l -5,5 v 15212 l 5,-6343 v 6348 l -5,-5 H 459 l 4896,5 H 454 l 5,-5 V 1791 l -5,7145 V 1787 h 1"
         id="path4118" />
    </clipPath>
    <mask
       maskUnits="userSpaceOnUse"
       x="0"
       y="0"
       width="1"
       height="1"
       id="mask4124">
      <image
         width="1"
         height="1"
         style="image-rendering:optimizeSpeed"
         preserveAspectRatio="none"
         xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAADMAAAAzCAAAAAAfym/2AAAAAXNCSVQI5gpbmQAAAK5JREFUSIntls0OwyAMg+28/zuzw6oSZv7MpGmHcmhJ5Q8nSCUQMkobUgTypYhENB9xh1BVjgaA6NJ8hjTKOlsgSRrbSB2xlsiqtFyYntuJEbByuxcPy6aaWQiBsF3sei4r14ZHPj5TEPYOADxgflPPwzzMMcP//re1X64Zc7zPRNuIgHWSElduppNZD5PFQZ/bhNi8diDt9cY+fHcPmVOD+86Y4jTsYSLplV4Wghfl7RxRskCApwAAAABJRU5ErkJggg=="
         id="image4126" />
    </mask>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath8328">
      <path
         d="M 0,0 H 12727 V 19455 H 0 V 0"
         id="path8326" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath13088">
      <path
         d="M 0,0 H 12727 V 19455 H 0 V 0"
         id="path13086" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath13096">
      <path
         d="M 0,0 H 12727 V 19455 H 0 V 0"
         id="path13094" />
    </clipPath>
    <mask
       maskUnits="userSpaceOnUse"
       x="0"
       y="0"
       width="1"
       height="1"
       id="mask13100">
      <image
         width="1"
         height="1"
         style="image-rendering:optimizeSpeed"
         preserveAspectRatio="none"
         xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAACkAAAApCAAAAACNC18qAAAAAXNCSVQI5gpbmQAAAIFJREFUOI3t1cEKwCAMA9BkPz765ztMHSvVpjBv8+LBR0WskXDjbLP5BYYs0pw7Z7lyL8sEPpQZHJQp7JQ5bJQCvOmRoTGolAQMoAQBK+0ulQRsQ01QhYUT/fJbqd+mXLPUSzt6vvDitrz3QtoUEmxlfX4WMjm2Yc4HdPp3OOt+pAtM+xg4AWFDfwAAAABJRU5ErkJggg=="
         id="image13102" />
    </mask>
  </defs>
  <sodipodi:namedview
     id="namedview2342"
     pagecolor="#ffffff"
     bordercolor="#000000"
     borderopacity="0.25"
     inkscape:showpageshadow="2"
     inkscape:pageopacity="0.0"
     inkscape:pagecheckerboard="0"
     inkscape:deskcolor="#d1d1d1"
     showgrid="false"
     inkscape:zoom="0.50796569"
     inkscape:cx="472.47286"
     inkscape:cy="694.92883"
     inkscape:window-width="1920"
     inkscape:window-height="1009"
     inkscape:window-x="1912"
     inkscape:window-y="-8"
     inkscape:window-maximized="1"
     inkscape:current-layer="g2346" />
  <g
     id="g2346"
     inkscape:groupmode="layer"
     inkscape:label="5630 La Jolla Blvd"
     transform="matrix(0.08,0,0,-0.08,18.666666,1594.6667)">
    <g
       id="g2348">
      <g
         id="g2350"
         clip-path="url(#clipPath2354)">
        <path
           d="m 12203,8904 -421,802"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2356" />
        <path
           d="m 11608,10038 -175,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2358" />
        <path
           d="m 11259,10702 -175,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2360" />
        <path
           d="m 10910,11366 -872,1660"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2362" />
        <path
           d="m 9864,13358 -175,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2364" />
        <path
           d="m 9515,14022 -175,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2366" />
        <path
           d="m 9166,14686 -872,1660"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2368" />
        <path
           d="m 8120,16678 -175,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2370" />
        <path
           d="m 7771,17342 -175,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2372" />
        <path
           d="m 7422,18006 -487,927"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2374" />
        <path
           d="M 10224,1787 1216,18933"
           style="fill:none;stroke:#0000ff;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2376" />
        <path
           d="m 6835,1787 -39,73"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2378" />
        <path
           d="m 6622,2192 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2380" />
        <path
           d="m 6273,2856 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2382" />
        <path
           d="M 5924,3520 5052,5180"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2384" />
        <path
           d="m 4878,5512 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2386" />
        <path
           d="m 4529,6176 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2388" />
        <path
           d="M 4180,6840 3308,8500"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2390" />
        <path
           d="m 3134,8832 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2392" />
        <path
           d="m 2785,9496 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2394" />
        <path
           d="m 2436,10160 -872,1660"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2396" />
        <path
           d="m 1390,12152 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2398" />
        <path
           d="m 1041,12816 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2400" />
        <path
           d="m 692,13480 -238,454"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2402" />
        <path
           d="M 12203,8823 6893,18933"
           style="fill:none;stroke:#0000ff;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2404" />
        <path
           d="m 12157,2328 -174,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2406" />
        <path
           d="m 11808,2992 -872,1660"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2408" />
        <path
           d="m 10762,4984 -175,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2410" />
        <path
           d="m 10413,5648 -174,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2412" />
        <path
           d="M 10064,6312 9192,7972"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2414" />
        <path
           d="m 9018,8304 -174,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2416" />
        <path
           d="m 8669,8968 -174,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2418" />
        <path
           d="m 8320,9632 -872,1660"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2420" />
        <path
           d="m 7274,11624 -174,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2422" />
        <path
           d="m 6925,12288 -174,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2424" />
        <path
           d="m 6576,12951 -872,1660"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2426" />
        <path
           d="m 5530,14943 -174,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2428" />
        <path
           d="m 5181,15607 -174,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2430" />
        <path
           d="m 4832,16271 -872,1660"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2432" />
        <path
           d="m 3786,18263 -174,332"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2434" />
        <path
           d="m 3437,18927 -3,6"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2436" />
        <path
           d="M 12203,12049 8587,18933"
           style="fill:none;stroke:#0000ff;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2438" />
        <path
           d="m 12203,13662 -158,302"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2440" />
        <path
           d="m 11870,14296 -174,332"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2442" />
        <path
           d="m 11522,14960 -175,332"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2444" />
        <path
           d="m 11173,15624 -872,1660"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2446" />
        <path
           d="m 10126,17616 -174,332"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2448" />
        <path
           d="m 9778,18280 -175,332"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2450" />
        <path
           d="m 12165,18896 -20,37"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2452" />
        <path
           d="m 12203,8823 -13,25"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2454" />
        <path
           d="m 12016,9180 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2456" />
        <path
           d="m 11667,9844 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2458" />
        <path
           d="m 11318,10508 -872,1660"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2460" />
        <path
           d="m 10272,12500 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2462" />
        <path
           d="m 9923,13164 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2464" />
        <path
           d="m 9574,13828 -872,1660"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2466" />
        <path
           d="m 8528,15820 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2468" />
        <path
           d="m 8179,16484 -174,332"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2470" />
        <path
           d="m 7830,17148 -872,1660"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2472" />
        <path
           d="M 1470,18933 10478,1787"
           style="fill:none;stroke:#0000ff;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2474" />
        <path
           d="m 9207,1787 -80,152 -290,-152"
           style="fill:none;stroke:#0000ff;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2476" />
        <path
           d="m 8750,1787 217,113 -244,465 -266,-139 231,-439"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2478" />
        <path
           d="m 9729,1787 v 0"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2480" />
        <path
           d="m 9729,1787 -32,17 -34,14 -35,10 -37,6 -36,1 -37,-2 -36,-7 13,23 10,24 6,25 3,27 -2,26 -4,25 -9,25 -12,23 -15,22 -18,19 -21,16 -23,13 -24,9 -26,6 -26,3"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2482" />
        <path
           d="m 9334.8945,2111.7761 c -44.9756,157.115 -203.1005,253.324 -363.3066,221.0496 -160.207,-32.2744 -268.7461,-182.2044 -249.3789,-344.4782"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2484" />
        <path
           d="m 8722,1988 -26,16 -29,13 -30,9 -30,6 -31,2 -31,-2 -31,-6 -30,-9 -28,-13 -27,-17 -24,-19 -22,-22 -19,-25 -16,-27 -12,-28 -9,-30 -6,-31 -1,-18"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2486" />
        <path
           d="m 7388,5976 299,156 -105,200 -299,-157 105,-199"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2488" />
        <path
           d="m 6281,6066 531,279 -279,531 -531,-279 279,-531"
           style="fill:none;stroke:#0000ff;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2490" />
        <path
           d="m 5815.5698,6520.7344 c -89.2593,-44.3091 -135.9941,-144.4732 -112.6064,-241.3418 23.3877,-96.8682 110.6767,-164.6739 210.3203,-163.3745"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2492" />
        <path
           d="m 5913.5127,6115.9302 c -52.9902,-96.6709 -27.5772,-217.541 59.8555,-284.688 87.4326,-67.1475 210.7666,-60.5132 290.4921,15.625"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2494" />
        <path
           d="m 6262.7812,5847.144 c 25.8389,-98.0722 119.3614,-162.6289 220.2237,-152.0156 100.8623,10.6128 178.8994,93.2217 183.7593,194.5244"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2496" />
        <path
           d="m 6667.3071,5889.7192 c 68.1529,-55.8115 167.1197,-52.4536 231.333,7.8487 64.2134,60.3027 73.7754,158.8637 22.3511,230.3847"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2498" />
        <path
           d="m 6921.5019,6129.0059 c 128.9273,-17.6993 255.9087,43.5795 322.2725,155.5229 66.3643,111.9434 59.1895,252.7544 -18.209,357.3726 -77.3984,104.6181 -209.9507,152.6728 -336.4111,121.9609"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2500" />
        <path
           d="m 6889.0669,6764.3696 c 37.9609,55.4219 42.4062,127.2173 11.5723,186.8989 -30.8345,59.6817 -91.9629,97.5992 -159.1299,98.7066"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2502" />
        <path
           d="m 6741.8945,7049.7764 c -44.9751,157.1147 -203.1001,253.3237 -363.3066,221.0493 -160.207,-32.2744 -268.7461,-182.2046 -249.3789,-344.478"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2504" />
        <path
           d="m 6129.4204,6926.4492 c -112.2461,77.6441 -265.6362,53.7925 -349.0059,-54.269 -83.3691,-108.0616 -67.5166,-262.4839 36.0689,-351.3535"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2506" />
        <path
           d="m 6485,6470.5 c 0,30.6519 -24.8481,55.5 -55.5,55.5 -30.6519,0 -55.5,-24.8481 -55.5,-55.5 0,-30.6519 24.8481,-55.5 55.5,-55.5 30.6519,0 55.5,24.8481 55.5,55.5"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path2508" />
        <path
           d="m 6932,3214 -45,92"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2510" />
        <path
           d="m 6885,3310 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2512" />
        <path
           d="m 6801,3483 -76,156"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2514" />
        <path
           d="m 6433,4237 -51,105"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2516" />
        <path
           d="m 6380,4346 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2518" />
        <path
           d="m 6296,4519 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2520" />
        <path
           d="m 6212,4691 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2522" />
        <path
           d="m 6128,4864 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2524" />
        <path
           d="m 6043,5036 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2526" />
        <path
           d="m 5959,5209 -25,52"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2528" />
        <path
           d="m 7321,2636 -53,109"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2530" />
        <path
           d="m 7266,2749 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2532" />
        <path
           d="m 7182,2921 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2534" />
        <path
           d="m 7098,3094 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2536" />
        <path
           d="m 7014,3266 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2538" />
        <path
           d="m 6929,3439 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2540" />
        <path
           d="m 6845,3611 -23,49"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2542" />
        <path
           d="m 6530,4258 -19,40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2544" />
        <path
           d="m 6509,4302 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2546" />
        <path
           d="m 6424,4474 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2548" />
        <path
           d="m 6340,4647 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2550" />
        <path
           d="m 6256,4819 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2552" />
        <path
           d="m 6172,4992 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2554" />
        <path
           d="m 6088,5165 -58,117"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2556" />
        <path
           d="m 7418,2657 -22,43"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2558" />
        <path
           d="m 7394,2704 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2560" />
        <path
           d="m 7310,2877 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2562" />
        <path
           d="m 7226,3050 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2564" />
        <path
           d="m 7142,3222 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2566" />
        <path
           d="m 7058,3395 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2568" />
        <path
           d="m 6974,3567 -56,114"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2570" />
        <path
           d="m 6626,4279 -71,147"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2572" />
        <path
           d="m 6553,4430 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2574" />
        <path
           d="m 6469,4603 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2576" />
        <path
           d="m 6384,4775 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2578" />
        <path
           d="m 6300,4948 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2580" />
        <path
           d="m 6216,5120 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2582" />
        <path
           d="m 6132,5293 -5,10"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2584" />
        <path
           d="m 7514,2678 -73,151"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2586" />
        <path
           d="m 7439,2833 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2588" />
        <path
           d="m 7354,3005 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2590" />
        <path
           d="m 7270,3178 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2592" />
        <path
           d="m 7186,3350 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2594" />
        <path
           d="m 7102,3523 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2596" />
        <path
           d="m 7018,3696 -3,6"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2598" />
        <path
           d="m 6723,4300 -40,82"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2600" />
        <path
           d="m 6681,4386 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2602" />
        <path
           d="m 6597,4558 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2604" />
        <path
           d="m 6513,4731 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2606" />
        <path
           d="m 6429,4904 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2608" />
        <path
           d="m 6344,5076 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2610" />
        <path
           d="m 6260,5249 -36,75"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2612" />
        <path
           d="m 7611,2699 -42,85"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2614" />
        <path
           d="m 7567,2789 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2616" />
        <path
           d="m 7483,2961 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2618" />
        <path
           d="m 7399,3134 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2620" />
        <path
           d="m 7315,3306 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2622" />
        <path
           d="m 7230,3479 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2624" />
        <path
           d="m 7146,3651 -35,72"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2626" />
        <path
           d="m 6820,4321 -9,17"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2628" />
        <path
           d="m 6809,4342 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2630" />
        <path
           d="m 6725,4514 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2632" />
        <path
           d="m 6641,4687 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2634" />
        <path
           d="m 6557,4859 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2636" />
        <path
           d="m 6473,5032 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2638" />
        <path
           d="m 6389,5205 -69,140"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2640" />
        <path
           d="m 7707,2720 -10,20"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2642" />
        <path
           d="m 7695,2744 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2644" />
        <path
           d="m 7611,2917 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2646" />
        <path
           d="m 7527,3089 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2648" />
        <path
           d="m 7443,3262 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2650" />
        <path
           d="m 7359,3435 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2652" />
        <path
           d="m 7275,3607 -67,137"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2654" />
        <path
           d="m 6916,4342 -60,124"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2656" />
        <path
           d="m 6854,4470 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2658" />
        <path
           d="m 6770,4643 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2660" />
        <path
           d="m 6685,4815 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2662" />
        <path
           d="m 6601,4988 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2664" />
        <path
           d="m 6517,5160 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2666" />
        <path
           d="m 6433,5333 -16,33"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2668" />
        <path
           d="m 7804,2741 -62,128"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2670" />
        <path
           d="m 7740,2873 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2672" />
        <path
           d="m 7655,3045 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2674" />
        <path
           d="m 7571,3218 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2676" />
        <path
           d="m 7487,3390 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2678" />
        <path
           d="m 7403,3563 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2680" />
        <path
           d="m 7319,3736 -15,29"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2682" />
        <path
           d="m 7013,4363 -29,59"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2684" />
        <path
           d="m 6982,4426 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2686" />
        <path
           d="m 6898,4598 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2688" />
        <path
           d="m 6814,4771 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2690" />
        <path
           d="m 6730,4944 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2692" />
        <path
           d="m 6645,5116 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2694" />
        <path
           d="m 6561,5289 -48,98"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2696" />
        <path
           d="m 7900,2762 -30,62"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2698" />
        <path
           d="m 7868,2829 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2700" />
        <path
           d="m 7784,3001 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2702" />
        <path
           d="m 7700,3174 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2704" />
        <path
           d="m 7615,3346 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2706" />
        <path
           d="m 7531,3519 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2708" />
        <path
           d="m 7447,3691 -46,95"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2710" />
        <path
           d="m 7109,4384 -81,166"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2712" />
        <path
           d="m 7026,4554 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2714" />
        <path
           d="m 6942,4727 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2716" />
        <path
           d="m 6858,4899 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2718" />
        <path
           d="m 6774,5072 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2720" />
        <path
           d="m 6690,5245 -80,163"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2722" />
        <path
           d="m 7996,2784 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2724" />
        <path
           d="m 7912,2957 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2726" />
        <path
           d="m 7828,3129 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2728" />
        <path
           d="m 7744,3302 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2730" />
        <path
           d="m 7660,3475 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2732" />
        <path
           d="m 7575,3647 -77,160"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2734" />
        <path
           d="m 7206,4405 -49,101"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2736" />
        <path
           d="m 7155,4510 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2738" />
        <path
           d="m 7070,4683 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2740" />
        <path
           d="m 6986,4855 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2742" />
        <path
           d="m 6902,5028 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2744" />
        <path
           d="m 6818,5200 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2746" />
        <path
           d="m 6734,5373 -28,56"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2748" />
        <path
           d="m 8094,2804 -51,105"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2750" />
        <path
           d="m 8041,2913 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2752" />
        <path
           d="m 7956,3085 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2754" />
        <path
           d="m 7872,3258 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2756" />
        <path
           d="m 7788,3430 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2758" />
        <path
           d="m 7704,3603 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2760" />
        <path
           d="m 7620,3776 -26,52"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2762" />
        <path
           d="m 7302,4426 -17,36"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2764" />
        <path
           d="m 7283,4466 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2766" />
        <path
           d="m 7199,4638 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2768" />
        <path
           d="m 7115,4811 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2770" />
        <path
           d="m 7030,4984 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2772" />
        <path
           d="m 6946,5156 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2774" />
        <path
           d="m 6862,5329 -59,121"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2776" />
        <path
           d="m 8190,2825 -19,39"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2778" />
        <path
           d="m 8169,2868 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2780" />
        <path
           d="m 8085,3041 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2782" />
        <path
           d="m 8001,3214 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2784" />
        <path
           d="m 7916,3386 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2786" />
        <path
           d="m 7832,3559 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2788" />
        <path
           d="m 7748,3731 -57,118"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2790" />
        <path
           d="m 7399,4447 -70,143"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2792" />
        <path
           d="m 7327,4594 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2794" />
        <path
           d="m 7243,4767 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2796" />
        <path
           d="m 7159,4939 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2798" />
        <path
           d="m 7075,5112 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2800" />
        <path
           d="m 6991,5285 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2802" />
        <path
           d="m 6906,5457 -6,14"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2804" />
        <path
           d="m 8287,2846 -72,147"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2806" />
        <path
           d="m 8213,2997 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2808" />
        <path
           d="m 8129,3169 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2810" />
        <path
           d="m 8045,3342 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2812" />
        <path
           d="m 7961,3515 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2814" />
        <path
           d="m 7876,3687 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2816" />
        <path
           d="m 7792,3860 -5,10"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2818" />
        <path
           d="m 7496,4468 -38,78"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2820" />
        <path
           d="m 7456,4550 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2822" />
        <path
           d="m 7371,4723 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2824" />
        <path
           d="m 7287,4895 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2826" />
        <path
           d="m 7203,5068 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2828" />
        <path
           d="m 7119,5240 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2830" />
        <path
           d="m 7035,5413 -39,79"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2832" />
        <path
           d="m 8383,2867 -40,82"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2834" />
        <path
           d="m 8341,2953 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2836" />
        <path
           d="m 8257,3125 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2838" />
        <path
           d="m 8173,3298 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2840" />
        <path
           d="m 8089,3470 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2842" />
        <path
           d="m 8005,3643 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2844" />
        <path
           d="m 7921,3816 -37,75"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2846" />
        <path
           d="m 7592,4489 -6,13"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2848" />
        <path
           d="m 7584,4506 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2850" />
        <path
           d="m 7500,4678 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2852" />
        <path
           d="m 7416,4851 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2854" />
        <path
           d="m 7331,5024 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2856" />
        <path
           d="m 7247,5196 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2858" />
        <path
           d="m 7163,5369 -70,144"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2860" />
        <path
           d="m 8480,2888 -8,16"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2862" />
        <path
           d="m 8470,2908 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2864" />
        <path
           d="m 8386,3081 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2866" />
        <path
           d="m 8302,3254 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2868" />
        <path
           d="m 8217,3426 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2870" />
        <path
           d="m 8133,3599 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2872" />
        <path
           d="m 8049,3771 -69,141"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2874" />
        <path
           d="m 7689,4510 -59,120"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2876" />
        <path
           d="m 7628,4634 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2878" />
        <path
           d="m 7544,4807 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2880" />
        <path
           d="m 7460,4979 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2882" />
        <path
           d="m 7376,5152 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2884" />
        <path
           d="m 7291,5324 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2886" />
        <path
           d="m 7207,5497 -18,37"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2888" />
        <path
           d="m 8577,2909 -61,124"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2890" />
        <path
           d="m 8514,3037 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2892" />
        <path
           d="m 8430,3209 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2894" />
        <path
           d="m 8346,3382 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2896" />
        <path
           d="m 8262,3555 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2898" />
        <path
           d="m 8177,3727 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2900" />
        <path
           d="m 8093,3900 -16,33"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2902" />
        <path
           d="m 6862,3347 -21,44"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2904" />
        <path
           d="m 6839,3395 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2906" />
        <path
           d="m 6755,3567 -35,71"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2908" />
        <path
           d="m 6429,4236 -9,18"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2910" />
        <path
           d="m 6418,4258 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2912" />
        <path
           d="m 6334,4430 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2914" />
        <path
           d="m 6250,4603 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2916" />
        <path
           d="m 6166,4775 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2918" />
        <path
           d="m 6082,4948 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2920" />
        <path
           d="m 5997,5121 -68,139"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2922" />
        <path
           d="m 7317,2635 -11,21"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2924" />
        <path
           d="m 7304,2660 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2926" />
        <path
           d="m 7220,2833 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2928" />
        <path
           d="m 7136,3005 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2930" />
        <path
           d="m 7052,3178 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2932" />
        <path
           d="m 6967,3351 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2934" />
        <path
           d="m 6883,3523 -66,136"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2936" />
        <path
           d="m 6525,4257 -61,125"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2938" />
        <path
           d="m 6462,4386 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2940" />
        <path
           d="m 6378,4559 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2942" />
        <path
           d="m 6294,4731 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2944" />
        <path
           d="m 6210,4904 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2946" />
        <path
           d="m 6126,5076 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2948" />
        <path
           d="m 6042,5249 -16,32"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2950" />
        <path
           d="m 7413,2656 -63,129"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2952" />
        <path
           d="m 7348,2789 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2954" />
        <path
           d="m 7264,2961 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2956" />
        <path
           d="m 7180,3134 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2958" />
        <path
           d="m 7096,3306 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2960" />
        <path
           d="m 7012,3479 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2962" />
        <path
           d="m 6927,3652 -13,28"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2964" />
        <path
           d="m 6622,4278 -29,60"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2966" />
        <path
           d="m 6591,4342 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2968" />
        <path
           d="m 6507,4514 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2970" />
        <path
           d="m 6422,4687 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2972" />
        <path
           d="m 6338,4860 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2974" />
        <path
           d="m 6254,5032 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2976" />
        <path
           d="m 6170,5205 -48,97"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2978" />
        <path
           d="m 7510,2677 -31,63"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2980" />
        <path
           d="m 7477,2744 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2982" />
        <path
           d="m 7393,2917 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2984" />
        <path
           d="m 7308,3090 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2986" />
        <path
           d="m 7224,3262 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2988" />
        <path
           d="m 7140,3435 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2990" />
        <path
           d="m 7056,3607 -46,94"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2992" />
        <path
           d="m 6718,4299 -81,167"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2994" />
        <path
           d="m 6635,4470 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2996" />
        <path
           d="m 6551,4643 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path2998" />
        <path
           d="m 6467,4815 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3000" />
        <path
           d="m 6382,4988 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3002" />
        <path
           d="m 6298,5161 -79,162"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3004" />
        <path
           d="m 7605,2700 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3006" />
        <path
           d="m 7521,2873 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3008" />
        <path
           d="m 7437,3045 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3010" />
        <path
           d="m 7353,3218 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3012" />
        <path
           d="m 7268,3391 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3014" />
        <path
           d="m 7184,3563 -77,159"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3016" />
        <path
           d="m 6815,4320 -50,102"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3018" />
        <path
           d="m 6763,4426 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3020" />
        <path
           d="m 6679,4599 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3022" />
        <path
           d="m 6595,4771 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3024" />
        <path
           d="m 6511,4944 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3026" />
        <path
           d="m 6427,5116 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3028" />
        <path
           d="m 6343,5289 -27,55"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3030" />
        <path
           d="m 7703,2719 -52,106"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3032" />
        <path
           d="m 7649,2829 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3034" />
        <path
           d="m 7565,3001 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3036" />
        <path
           d="m 7481,3174 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3038" />
        <path
           d="m 7397,3346 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3040" />
        <path
           d="m 7313,3519 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3042" />
        <path
           d="m 7228,3692 -25,51"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3044" />
        <path
           d="m 6912,4341 -18,37"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3046" />
        <path
           d="m 6892,4382 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3048" />
        <path
           d="m 6808,4554 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3050" />
        <path
           d="m 6723,4727 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3052" />
        <path
           d="m 6639,4900 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3054" />
        <path
           d="m 6555,5072 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3056" />
        <path
           d="m 6471,5245 -59,120"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3058" />
        <path
           d="m 7799,2740 -19,40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3060" />
        <path
           d="m 7778,2784 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3062" />
        <path
           d="m 7693,2957 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3064" />
        <path
           d="m 7609,3130 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3066" />
        <path
           d="m 7525,3302 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3068" />
        <path
           d="m 7441,3475 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3070" />
        <path
           d="m 7357,3647 -57,117"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3072" />
        <path
           d="m 7008,4362 -70,144"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3074" />
        <path
           d="m 6936,4510 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3076" />
        <path
           d="m 6852,4683 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3078" />
        <path
           d="m 6768,4855 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3080" />
        <path
           d="m 6683,5028 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3082" />
        <path
           d="m 6599,5200 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3084" />
        <path
           d="m 6515,5373 -6,13"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3086" />
        <path
           d="m 7896,2761 -72,148"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3088" />
        <path
           d="m 7822,2913 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3090" />
        <path
           d="m 7738,3085 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3092" />
        <path
           d="m 7653,3258 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3094" />
        <path
           d="m 7569,3431 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3096" />
        <path
           d="m 7485,3603 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3098" />
        <path
           d="m 7401,3776 -4,9"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3100" />
        <path
           d="m 7105,4383 -39,79"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3102" />
        <path
           d="m 7064,4466 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3104" />
        <path
           d="m 6980,4639 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3106" />
        <path
           d="m 6896,4811 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3108" />
        <path
           d="m 6812,4984 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3110" />
        <path
           d="m 6728,5156 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3112" />
        <path
           d="m 6643,5329 -38,78"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3114" />
        <path
           d="m 7993,2782 -41,83"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3116" />
        <path
           d="m 7950,2869 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3118" />
        <path
           d="m 7866,3041 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3120" />
        <path
           d="m 7782,3214 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3122" />
        <path
           d="m 7698,3386 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3124" />
        <path
           d="m 7614,3559 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3126" />
        <path
           d="m 7529,3731 -36,75"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3128" />
        <path
           d="m 7201,4404 -6,14"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3130" />
        <path
           d="m 7193,4422 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3132" />
        <path
           d="m 7109,4594 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3134" />
        <path
           d="m 7024,4767 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3136" />
        <path
           d="m 6940,4940 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3138" />
        <path
           d="m 6856,5112 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3140" />
        <path
           d="m 6772,5285 -70,143"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3142" />
        <path
           d="m 8089,2803 -8,17"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3144" />
        <path
           d="m 8079,2824 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3146" />
        <path
           d="m 7994,2997 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3148" />
        <path
           d="m 7910,3170 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3150" />
        <path
           d="m 7826,3342 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3152" />
        <path
           d="m 7742,3515 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3154" />
        <path
           d="m 7658,3687 -68,140"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3156" />
        <path
           d="m 7298,4425 -59,121"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3158" />
        <path
           d="m 7237,4550 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3160" />
        <path
           d="m 7153,4723 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3162" />
        <path
           d="m 7069,4895 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3164" />
        <path
           d="m 6984,5068 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3166" />
        <path
           d="m 6900,5240 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3168" />
        <path
           d="m 6816,5413 -18,36"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3170" />
        <path
           d="m 8186,2824 -61,125"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3172" />
        <path
           d="m 8123,2953 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3174" />
        <path
           d="m 8039,3125 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3176" />
        <path
           d="m 7954,3298 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3178" />
        <path
           d="m 7870,3471 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3180" />
        <path
           d="m 7786,3643 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3182" />
        <path
           d="m 7702,3816 -16,32"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3184" />
        <path
           d="m 7395,4446 -28,56"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3186" />
        <path
           d="m 7365,4506 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3188" />
        <path
           d="m 7281,4679 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3190" />
        <path
           d="m 7197,4851 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3192" />
        <path
           d="m 7113,5024 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3194" />
        <path
           d="m 7029,5196 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3196" />
        <path
           d="m 6944,5369 -49,101"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3198" />
        <path
           d="m 8282,2845 -29,60"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3200" />
        <path
           d="m 8251,2909 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3202" />
        <path
           d="m 8167,3081 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3204" />
        <path
           d="m 8083,3254 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3206" />
        <path
           d="m 7999,3426 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3208" />
        <path
           d="m 7914,3599 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3210" />
        <path
           d="m 7830,3771 -47,98"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3212" />
        <path
           d="m 7491,4467 -80,163"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3214" />
        <path
           d="m 7409,4634 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3216" />
        <path
           d="m 7325,4807 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3218" />
        <path
           d="m 7241,4979 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3220" />
        <path
           d="m 7157,5152 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3222" />
        <path
           d="m 7073,5325 -81,166"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3224" />
        <path
           d="m 8379,2866 -82,167"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3226" />
        <path
           d="m 8295,3037 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3228" />
        <path
           d="m 8211,3210 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3230" />
        <path
           d="m 8127,3382 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3232" />
        <path
           d="m 8043,3555 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3234" />
        <path
           d="m 7959,3727 -80,163"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3236" />
        <path
           d="m 7588,4488 -48,98"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3238" />
        <path
           d="m 7538,4590 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3240" />
        <path
           d="m 7454,4763 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3242" />
        <path
           d="m 7369,4935 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3244" />
        <path
           d="m 7285,5108 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3246" />
        <path
           d="m 7201,5280 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3248" />
        <path
           d="m 7117,5453 -29,59"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3250" />
        <path
           d="m 8475,2887 -49,102"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3252" />
        <path
           d="m 8424,2993 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3254" />
        <path
           d="m 8340,3165 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3256" />
        <path
           d="m 8255,3338 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3258" />
        <path
           d="m 8171,3510 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3260" />
        <path
           d="m 8087,3683 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3262" />
        <path
           d="m 8003,3856 -27,55"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3264" />
        <path
           d="m 7684,4509 -16,33"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3266" />
        <path
           d="m 7666,4546 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3268" />
        <path
           d="m 7582,4718 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3270" />
        <path
           d="m 7498,4891 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3272" />
        <path
           d="m 7414,5064 -83,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3274" />
        <path
           d="m 7330,5236 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3276" />
        <path
           d="m 7245,5409 -60,124"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3278" />
        <path
           d="m 8572,2908 -18,37"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3280" />
        <path
           d="m 8552,2949 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3282" />
        <path
           d="m 8468,3121 -82,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3284" />
        <path
           d="m 8384,3294 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3286" />
        <path
           d="m 8300,3466 -83,169"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3288" />
        <path
           d="m 8215,3639 -82,168"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3290" />
        <path
           d="m 8131,3811 -58,121"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3292" />
        <path
           d="m 8552,2949 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3294" />
        <path
           d="m 8543,3051 -29,-14"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3296" />
        <path
           d="m 8424,2993 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3298" />
        <path
           d="m 8251,2909 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3300" />
        <path
           d="m 8079,2824 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3302" />
        <path
           d="m 8468,3121 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3304" />
        <path
           d="m 8295,3037 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3306" />
        <path
           d="m 8123,2953 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3308" />
        <path
           d="m 7950,2869 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3310" />
        <path
           d="m 7778,2784 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3312" />
        <path
           d="m 7605,2700 -10,-5"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3314" />
        <path
           d="m 8454,3221 -24,-12"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3316" />
        <path
           d="m 8340,3165 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3318" />
        <path
           d="m 8167,3081 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3320" />
        <path
           d="m 7994,2997 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3322" />
        <path
           d="m 7822,2913 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3324" />
        <path
           d="m 7649,2829 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3326" />
        <path
           d="m 7477,2744 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3328" />
        <path
           d="m 7304,2660 -64,-31"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3330" />
        <path
           d="m 8384,3294 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3332" />
        <path
           d="m 8211,3210 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3334" />
        <path
           d="m 8039,3125 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3336" />
        <path
           d="m 7866,3041 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3338" />
        <path
           d="m 7693,2957 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3340" />
        <path
           d="m 7521,2873 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3342" />
        <path
           d="m 7348,2789 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3344" />
        <path
           d="m 8364,3391 -18,-9"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3346" />
        <path
           d="m 8255,3338 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3348" />
        <path
           d="m 8083,3254 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3350" />
        <path
           d="m 7910,3170 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3352" />
        <path
           d="m 7738,3085 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3354" />
        <path
           d="m 7565,3001 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3356" />
        <path
           d="m 7393,2917 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3358" />
        <path
           d="m 7220,2833 -70,-34"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3360" />
        <path
           d="m 8300,3466 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3362" />
        <path
           d="m 8127,3382 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3364" />
        <path
           d="m 7954,3298 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3366" />
        <path
           d="m 7782,3214 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3368" />
        <path
           d="m 7609,3130 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3370" />
        <path
           d="m 7437,3045 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3372" />
        <path
           d="m 7264,2961 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3374" />
        <path
           d="m 8275,3561 -13,-6"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3376" />
        <path
           d="m 8171,3510 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3378" />
        <path
           d="m 7999,3426 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3380" />
        <path
           d="m 7826,3342 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3382" />
        <path
           d="m 7653,3258 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3384" />
        <path
           d="m 7481,3174 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3386" />
        <path
           d="m 7308,3090 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3388" />
        <path
           d="m 7136,3005 -75,-36"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3390" />
        <path
           d="m 8215,3639 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3392" />
        <path
           d="m 8043,3555 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3394" />
        <path
           d="m 7870,3471 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3396" />
        <path
           d="m 7698,3386 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3398" />
        <path
           d="m 7525,3302 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3400" />
        <path
           d="m 7353,3218 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3402" />
        <path
           d="m 7180,3134 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3404" />
        <path
           d="m 8186,3731 -9,-4"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3406" />
        <path
           d="m 8087,3683 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3408" />
        <path
           d="m 7914,3599 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3410" />
        <path
           d="m 7742,3515 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3412" />
        <path
           d="m 7569,3431 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3414" />
        <path
           d="m 7397,3346 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3416" />
        <path
           d="m 7224,3262 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3418" />
        <path
           d="m 7052,3178 -80,-39"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3420" />
        <path
           d="m 8131,3811 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3422" />
        <path
           d="m 7959,3727 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3424" />
        <path
           d="m 7786,3643 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3426" />
        <path
           d="m 7614,3559 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3428" />
        <path
           d="m 7441,3475 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3430" />
        <path
           d="m 7268,3391 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3432" />
        <path
           d="m 7096,3306 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3434" />
        <path
           d="m 8096,3901 -3,-1"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3436" />
        <path
           d="m 8003,3856 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3438" />
        <path
           d="m 7830,3771 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3440" />
        <path
           d="m 7658,3687 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3442" />
        <path
           d="m 7485,3603 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3444" />
        <path
           d="m 7313,3519 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3446" />
        <path
           d="m 7140,3435 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3448" />
        <path
           d="m 6967,3351 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3450" />
        <path
           d="m 7834,3880 -42,-20"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3452" />
        <path
           d="m 7702,3816 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3454" />
        <path
           d="m 7529,3731 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3456" />
        <path
           d="m 7357,3647 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3458" />
        <path
           d="m 7184,3563 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3460" />
        <path
           d="m 7012,3479 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3462" />
        <path
           d="m 6839,3395 -1,-1"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3464" />
        <path
           d="m 7401,3776 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3466" />
        <path
           d="m 7228,3692 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3468" />
        <path
           d="m 7056,3607 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3470" />
        <path
           d="m 6883,3523 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3472" />
        <path
           d="m 7044,3708 -26,-12"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3474" />
        <path
           d="m 6927,3652 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3476" />
        <path
           d="m 6755,3567 -7,-3"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3478" />
        <path
           d="m 7666,4546 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3480" />
        <path
           d="m 7694,4666 -66,-32"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3482" />
        <path
           d="m 7538,4590 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3484" />
        <path
           d="m 7365,4506 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3486" />
        <path
           d="m 7193,4422 -73,-36"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3488" />
        <path
           d="m 7582,4718 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3490" />
        <path
           d="m 7409,4634 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3492" />
        <path
           d="m 7237,4550 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3494" />
        <path
           d="m 7064,4466 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3496" />
        <path
           d="m 6892,4382 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3498" />
        <path
           d="m 7605,4836 -61,-29"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3500" />
        <path
           d="m 7454,4763 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3502" />
        <path
           d="m 7281,4679 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3504" />
        <path
           d="m 7109,4594 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3506" />
        <path
           d="m 6936,4510 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3508" />
        <path
           d="m 6763,4426 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3510" />
        <path
           d="m 6591,4342 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3512" />
        <path
           d="m 6418,4258 -27,-14"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3514" />
        <path
           d="m 7498,4891 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3516" />
        <path
           d="m 7325,4807 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3518" />
        <path
           d="m 7153,4723 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3520" />
        <path
           d="m 6980,4639 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3522" />
        <path
           d="m 6808,4554 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3524" />
        <path
           d="m 6635,4470 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3526" />
        <path
           d="m 6462,4386 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3528" />
        <path
           d="m 7516,5007 -56,-28"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3530" />
        <path
           d="m 7369,4935 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3532" />
        <path
           d="m 7197,4851 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3534" />
        <path
           d="m 7024,4767 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3536" />
        <path
           d="m 6852,4683 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3538" />
        <path
           d="m 6679,4599 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3540" />
        <path
           d="m 6507,4514 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3542" />
        <path
           d="m 6334,4430 -32,-16"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3544" />
        <path
           d="m 7414,5064 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3546" />
        <path
           d="m 7241,4979 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3548" />
        <path
           d="m 7069,4895 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3550" />
        <path
           d="m 6896,4811 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3552" />
        <path
           d="m 6723,4727 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3554" />
        <path
           d="m 6551,4643 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3556" />
        <path
           d="m 6378,4559 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3558" />
        <path
           d="m 7426,5177 -50,-25"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3560" />
        <path
           d="m 7285,5108 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3562" />
        <path
           d="m 7113,5024 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3564" />
        <path
           d="m 6940,4940 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3566" />
        <path
           d="m 6768,4855 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3568" />
        <path
           d="m 6595,4771 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3570" />
        <path
           d="m 6422,4687 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3572" />
        <path
           d="m 6250,4603 -38,-18"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3574" />
        <path
           d="m 7330,5236 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3576" />
        <path
           d="m 7157,5152 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3578" />
        <path
           d="m 6984,5068 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3580" />
        <path
           d="m 6812,4984 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3582" />
        <path
           d="m 6639,4900 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3584" />
        <path
           d="m 6467,4815 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3586" />
        <path
           d="m 6294,4731 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3588" />
        <path
           d="m 7337,5347 -46,-23"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3590" />
        <path
           d="m 7201,5280 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3592" />
        <path
           d="m 7029,5196 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3594" />
        <path
           d="m 6856,5112 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3596" />
        <path
           d="m 6683,5028 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3598" />
        <path
           d="m 6511,4944 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3600" />
        <path
           d="m 6338,4860 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3602" />
        <path
           d="m 6166,4775 -43,-20"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3604" />
        <path
           d="m 7245,5409 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3606" />
        <path
           d="m 7073,5325 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3608" />
        <path
           d="m 6900,5240 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3610" />
        <path
           d="m 6728,5156 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3612" />
        <path
           d="m 6555,5072 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3614" />
        <path
           d="m 6382,4988 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3616" />
        <path
           d="m 6210,4904 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3618" />
        <path
           d="m 7248,5517 -41,-20"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3620" />
        <path
           d="m 7117,5453 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3622" />
        <path
           d="m 6944,5369 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3624" />
        <path
           d="m 6772,5285 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3626" />
        <path
           d="m 6599,5200 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3628" />
        <path
           d="m 6427,5116 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3630" />
        <path
           d="m 6254,5032 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3632" />
        <path
           d="m 6082,4948 -48,-23"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3634" />
        <path
           d="m 6963,5485 -57,-28"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3636" />
        <path
           d="m 6816,5413 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3638" />
        <path
           d="m 6643,5329 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3640" />
        <path
           d="m 6471,5245 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3642" />
        <path
           d="m 6298,5161 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3644" />
        <path
           d="m 6126,5076 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3646" />
        <path
           d="m 6515,5373 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3648" />
        <path
           d="m 6343,5289 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3650" />
        <path
           d="m 6170,5205 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3652" />
        <path
           d="m 5997,5121 -53,-26"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3654" />
        <path
           d="m 6173,5313 -41,-20"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3656" />
        <path
           d="m 6042,5249 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3658" />
        <path
           d="m 8554,2945 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3660" />
        <path
           d="m 8545,3047 -29,-14"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3662" />
        <path
           d="m 8426,2989 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3664" />
        <path
           d="m 8253,2905 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3666" />
        <path
           d="m 8081,2820 -72,-35"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3668" />
        <path
           d="m 8470,3117 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3670" />
        <path
           d="m 8297,3033 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3672" />
        <path
           d="m 8125,2949 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3674" />
        <path
           d="m 7952,2865 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3676" />
        <path
           d="m 7780,2780 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3678" />
        <path
           d="m 8456,3217 -24,-12"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3680" />
        <path
           d="m 8342,3161 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3682" />
        <path
           d="m 8169,3077 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3684" />
        <path
           d="m 7996,2993 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3686" />
        <path
           d="m 7824,2909 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3688" />
        <path
           d="m 7651,2825 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3690" />
        <path
           d="m 7479,2740 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3692" />
        <path
           d="m 7306,2656 -64,-31"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3694" />
        <path
           d="m 8386,3290 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3696" />
        <path
           d="m 8213,3205 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3698" />
        <path
           d="m 8041,3121 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3700" />
        <path
           d="m 7868,3037 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3702" />
        <path
           d="m 7695,2953 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3704" />
        <path
           d="m 7523,2869 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3706" />
        <path
           d="m 7350,2785 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3708" />
        <path
           d="m 8366,3387 -18,-9"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3710" />
        <path
           d="m 8257,3334 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3712" />
        <path
           d="m 8085,3250 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3714" />
        <path
           d="m 7912,3166 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3716" />
        <path
           d="m 7740,3081 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3718" />
        <path
           d="m 7567,2997 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3720" />
        <path
           d="m 7394,2913 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3722" />
        <path
           d="m 7222,2829 -70,-34"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3724" />
        <path
           d="m 8302,3462 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3726" />
        <path
           d="m 8129,3378 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3728" />
        <path
           d="m 7956,3294 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3730" />
        <path
           d="m 7784,3210 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3732" />
        <path
           d="m 7611,3126 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3734" />
        <path
           d="m 7439,3041 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3736" />
        <path
           d="m 7266,2957 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3738" />
        <path
           d="m 8277,3557 -13,-7"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3740" />
        <path
           d="m 8173,3506 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3742" />
        <path
           d="m 8001,3422 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3744" />
        <path
           d="m 7828,3338 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3746" />
        <path
           d="m 7655,3254 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3748" />
        <path
           d="m 7483,3170 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3750" />
        <path
           d="m 7310,3086 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3752" />
        <path
           d="m 7138,3001 -75,-36"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3754" />
        <path
           d="m 8217,3635 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3756" />
        <path
           d="m 8045,3551 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3758" />
        <path
           d="m 7872,3466 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3760" />
        <path
           d="m 7700,3382 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3762" />
        <path
           d="m 7527,3298 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3764" />
        <path
           d="m 7355,3214 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3766" />
        <path
           d="m 7182,3130 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3768" />
        <path
           d="m 8188,3727 -9,-4"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3770" />
        <path
           d="m 8089,3679 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3772" />
        <path
           d="m 7916,3595 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3774" />
        <path
           d="m 7744,3511 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3776" />
        <path
           d="m 7571,3427 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3778" />
        <path
           d="m 7399,3342 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3780" />
        <path
           d="m 7226,3258 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3782" />
        <path
           d="m 7054,3174 -80,-39"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3784" />
        <path
           d="m 8133,3807 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3786" />
        <path
           d="m 7961,3723 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3788" />
        <path
           d="m 7788,3639 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3790" />
        <path
           d="m 7615,3555 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3792" />
        <path
           d="m 7443,3471 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3794" />
        <path
           d="m 7270,3387 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3796" />
        <path
           d="m 7098,3302 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3798" />
        <path
           d="m 8098,3897 -3,-1"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3800" />
        <path
           d="m 8005,3852 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3802" />
        <path
           d="m 7832,3767 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3804" />
        <path
           d="m 7660,3683 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3806" />
        <path
           d="m 7487,3599 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3808" />
        <path
           d="m 7315,3515 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3810" />
        <path
           d="m 7142,3431 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3812" />
        <path
           d="m 6969,3347 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3814" />
        <path
           d="m 7852,3884 -58,-28"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3816" />
        <path
           d="m 7704,3812 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3818" />
        <path
           d="m 7531,3727 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3820" />
        <path
           d="m 7359,3643 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3822" />
        <path
           d="m 7186,3559 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3824" />
        <path
           d="m 7014,3475 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3826" />
        <path
           d="m 6841,3391 -1,-1"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3828" />
        <path
           d="m 7403,3772 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3830" />
        <path
           d="m 7230,3687 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3832" />
        <path
           d="m 7058,3603 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3834" />
        <path
           d="m 6885,3519 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3836" />
        <path
           d="m 7062,3712 -42,-20"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3838" />
        <path
           d="m 6929,3648 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3840" />
        <path
           d="m 6757,3563 -7,-3"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3842" />
        <path
           d="m 7668,4542 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3844" />
        <path
           d="m 7696,4662 -66,-32"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3846" />
        <path
           d="m 7540,4586 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3848" />
        <path
           d="m 7367,4502 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3850" />
        <path
           d="m 7195,4418 -57,-28"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3852" />
        <path
           d="m 7584,4714 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3854" />
        <path
           d="m 7411,4630 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3856" />
        <path
           d="m 7239,4546 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3858" />
        <path
           d="m 7066,4462 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3860" />
        <path
           d="m 6894,4378 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3862" />
        <path
           d="m 7607,4832 -61,-29"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3864" />
        <path
           d="m 7456,4759 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3866" />
        <path
           d="m 7283,4674 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3868" />
        <path
           d="m 7110,4590 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3870" />
        <path
           d="m 6938,4506 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3872" />
        <path
           d="m 6765,4422 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3874" />
        <path
           d="m 6593,4338 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3876" />
        <path
           d="m 6420,4254 -27,-14"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3878" />
        <path
           d="m 7500,4887 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3880" />
        <path
           d="m 7327,4803 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3882" />
        <path
           d="m 7155,4719 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3884" />
        <path
           d="m 6982,4635 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3886" />
        <path
           d="m 6810,4550 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3888" />
        <path
           d="m 6637,4466 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3890" />
        <path
           d="m 6464,4382 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3892" />
        <path
           d="m 7518,5003 -56,-28"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3894" />
        <path
           d="m 7371,4931 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3896" />
        <path
           d="m 7199,4847 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3898" />
        <path
           d="m 7026,4763 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3900" />
        <path
           d="m 6854,4679 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3902" />
        <path
           d="m 6681,4595 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3904" />
        <path
           d="m 6509,4510 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3906" />
        <path
           d="m 6336,4426 -32,-16"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3908" />
        <path
           d="m 7416,5060 -83,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3910" />
        <path
           d="m 7243,4975 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3912" />
        <path
           d="m 7071,4891 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3914" />
        <path
           d="m 6898,4807 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3916" />
        <path
           d="m 6725,4723 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3918" />
        <path
           d="m 6553,4639 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3920" />
        <path
           d="m 6380,4555 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3922" />
        <path
           d="m 7428,5173 -50,-25"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3924" />
        <path
           d="m 7287,5104 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3926" />
        <path
           d="m 7115,5020 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3928" />
        <path
           d="m 6942,4935 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3930" />
        <path
           d="m 6770,4851 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3932" />
        <path
           d="m 6597,4767 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3934" />
        <path
           d="m 6424,4683 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3936" />
        <path
           d="m 6252,4599 -38,-18"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3938" />
        <path
           d="m 7331,5232 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3940" />
        <path
           d="m 7159,5148 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3942" />
        <path
           d="m 6986,5064 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3944" />
        <path
           d="m 6814,4980 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3946" />
        <path
           d="m 6641,4895 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3948" />
        <path
           d="m 6469,4811 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3950" />
        <path
           d="m 6296,4727 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3952" />
        <path
           d="m 7339,5343 -46,-23"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3954" />
        <path
           d="m 7203,5276 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3956" />
        <path
           d="m 7031,5192 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3958" />
        <path
           d="m 6858,5108 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3960" />
        <path
           d="m 6685,5024 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3962" />
        <path
           d="m 6513,4940 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3964" />
        <path
           d="m 6340,4856 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3966" />
        <path
           d="m 6168,4771 -43,-20"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3968" />
        <path
           d="m 7247,5405 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3970" />
        <path
           d="m 7075,5321 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3972" />
        <path
           d="m 6902,5236 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3974" />
        <path
           d="m 6730,5152 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3976" />
        <path
           d="m 6557,5068 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3978" />
        <path
           d="m 6384,4984 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3980" />
        <path
           d="m 6212,4900 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3982" />
        <path
           d="m 7250,5513 -41,-20"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3984" />
        <path
           d="m 7119,5449 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3986" />
        <path
           d="m 6946,5365 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3988" />
        <path
           d="m 6774,5281 -82,-41"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3990" />
        <path
           d="m 6601,5196 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3992" />
        <path
           d="m 6429,5112 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3994" />
        <path
           d="m 6256,5028 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3996" />
        <path
           d="m 6084,4944 -48,-23"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path3998" />
        <path
           d="m 6982,5489 -74,-36"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4000" />
        <path
           d="m 6818,5409 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4002" />
        <path
           d="m 6645,5325 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4004" />
        <path
           d="m 6473,5241 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4006" />
        <path
           d="m 6300,5156 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4008" />
        <path
           d="m 6128,5072 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4010" />
        <path
           d="m 6517,5369 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4012" />
        <path
           d="m 6344,5285 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4014" />
        <path
           d="m 6172,5201 -82,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4016" />
        <path
           d="m 5999,5117 -53,-26"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4018" />
        <path
           d="m 6192,5317 -58,-28"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4020" />
        <path
           d="m 6044,5245 -83,-40"
           style="fill:none;stroke:#808080;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.24706"
           id="path4022" />
        <path
           d="M 7233,5544 7767,4527 6399,4230 5865,5246 7233,5544"
           style="fill:none;stroke:#0000ff;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4024" />
        <path
           d="M 8079,3933 6711,3636 7245,2619 8613,2917 8079,3933"
           style="fill:none;stroke:#0000ff;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4026" />
        <path
           d="M 9493,3177 9244,3046"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4028" />
        <path
           d="M 9078,2959 8746,2784"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4030" />
        <path
           d="M 8580,2697 8248,2523"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4032" />
        <path
           d="M 8082,2436 7751,2261"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4034" />
        <path
           d="M 7585,2174 7253,2000"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4036" />
        <path
           d="M 7087,1912 6847,1787"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4038" />
        <path
           d="M 9514,3137 9265,3006"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4040" />
        <path
           d="M 9099,2919 8767,2745"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4042" />
        <path
           d="M 8601,2657 8269,2483"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4044" />
        <path
           d="M 8103,2396 7771,2221"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4046" />
        <path
           d="M 7605,2134 7273,1960"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4048" />
        <path
           d="m 7107,1873 -163,-86"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4050" />
        <path
           d="M 9159,3814 8910,3683"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4052" />
        <path
           d="M 8744,3596 8412,3422"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4054" />
        <path
           d="M 8246,3334 7914,3160"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4056" />
        <path
           d="M 7748,3073 7416,2898"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4058" />
        <path
           d="M 7250,2811 6918,2637"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4060" />
        <path
           d="M 6752,2550 6503,2419"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4062" />
        <path
           d="M 9180,3774 8931,3643"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4064" />
        <path
           d="M 8765,3556 8433,3382"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4066" />
        <path
           d="M 8267,3294 7935,3120"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4068" />
        <path
           d="M 7769,3033 7437,2858"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4070" />
        <path
           d="M 7271,2771 6939,2597"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4072" />
        <path
           d="M 6773,2510 6524,2379"
           style="fill:none;stroke:#a500dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4074" />
      </g>
    </g>
    <g
       id="g4076">
      <g
         id="g4078"
         clip-path="url(#clipPath4082)" />
    </g>
    <g
       id="g4084">
      <g
         id="g4086"
         clip-path="url(#clipPath4090)">
        <g
           id="g4092"
           transform="matrix(153,0,0,153,7118,2928)">
          <image
             width="1"
             height="1"
             style="image-rendering:optimizeSpeed"
             preserveAspectRatio="none"
             transform="matrix(1,0,0,-1,0,1)"
             xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAADMAAAAzCAYAAAA6oTAqAAAABHNCSVQICAgIfAhkiAAADThJREFUaIGdWmtv28YSPeTyKZISJcuWH0lTow8gX/v/f0D/QFGgaJEgcGTZepiiRFHkkrv3gzpzVwyd5N4FBiJlmdyzM3PmsQsA+mvi+762LEsD0GEY8veDwYCvLy4uNABdFIWm0bat1lprpZRu25ZFKaXN0batdhzn7J2O4/A7XdfVAHSaphoAf9+9BqCtfy++OlzXhZQSAOB5HpqmgVIKjuOgLEs4joOXlxeMx2NorVEUBTzPw3w+x+Xl5dmzLMs6E9/3sd/vEccxwjDE8Xjkd2qt0TQNhBBo2xaWZSEIApRlCd/3UVXV+bO/BUYIAc/zUJYlwjCEUgpt22K73WIwGKBpGuR5jslkgvl8Dtd1oZRCkiRo2xZ1XX8BxrbtM0CO4yAMQwYVBAGqqjpbOAAYj8d4eXnh/9da89++C4w5qqpCXdeI4xi73Q5aawyHQ3z69AlhGCKKIhwOBwDAYrFAkiQQQkBrDcuyesEQ8CzLMJvN4LouDocDfN+H4zhn74/jGJ7nYbPZ9M7vm2BInVprZFmGNE2x3+9RVRUsy0JZlmjbFpvNBsPhEC8vL7i9vcV+v2dzM7XSBTMYDOD7PoqigO/78DwPQgg0TYM0Tfm3juOgaRoAQBiGbHamqX2XZo7HI3zfBwDM53NMJhOUZcma8n0feZ5DKYWyLKGUwnQ6xXq9ZjMwzcq2bZ4kAJRliZubG57wYDBAFEXIsgxN0+D29haO48CyLAaUpimyLPvfNEMOWNc1FosFLi4uUJYlNpsNHMdBXdc4HA4QQiAMQ0gp8fz8jDRNeSG6JmaCcV0Xw+EQy+USvu/j6uoK6/Ua9/f3aJoGQRBACMHPGA6HyPMcABBFEYqi+H4wWmtsNhskSYKqqrBer5lxtNZo2xa73Y41lGUZRqMRdrsdALDdd7VCYJRSiKIInuehKApEUYSrqys8Pj5iNpvBtm0kSQLgZPLEbPR5phkhhDbVNxgMYFkWPnz4gMvLS0gpUdc1yrJEXdeQUkJKiePxCCklmqZhIZPSWrNIKaH1f9fLBGPbNoQQcF0XrutCCMHs6fs+fN/HaDRCnueYzWZomgaHwwHT6RRCiDN/CYIAlmVZWmuN6+trLJdLtG3LprVareC6LqqqwvF4RFVVaJoGdV2zv9R1zWDatj0DopTiReqaGZkOsZbrunAch8EFQQDP82BZFqSUmE6nGAwGbMpELKPRCNvt9qRpnCIu2yeZVVVVUErxpE3NEBgpJYOna6UUA6GY1AVDGqBrx3GYxUgzBObi4oI1s9lsMBqNMJlM0LYtfN9nrQshwER+fX2NxWIBKSWyLEMcx2xKJgiaOAn5DWmGAJGQZshnKO5orWHb9plGSTNkjsApXk0mE+R5Dq01m91oNOIFCILgREie5zFTkY17nofj8Yj1es2M1iemzxBQUyNdMzO1YmqGtNm2LRMGEURZlphMJpBSIkkSbLdbCCFwPB6ZKSnmsGa01lgsFmyneZ7DdV0OkCRdn+kC62qma2ZdMLRYBMRxnDMiefPmDfuy53nwPA+73Q739/eYz+e4urrC8/PziQDwLzWT6pfLJRzHwePjI6/sawRgasb0GVNMJusSgG3baNsWruvC8zwG4/s+giCA7/uQUuLdu3eI4xhVVaFtW7x//x7r9RrT6RRPT0/47bffMJ/P4VAmejwe0TTNWbZK35MvdH2jaRr+OwEznZ/8oo+a27ZlU6Ln2bZ9ZqJKKQRBgCzLUJYlBoMBJpMJ/vnnH0wmExRFgdlshvl8fiIAskuiw6IosF6vcXl5idVqdZahUnwhQmiaBq0CZKNOIs/Z7PQpOXqfgOgzcRwHlgJaBVithoYCrBa2aKC0Bct2YDcKrmehaTW2+R5BEKBpNexGYblcciLrUEoihMBms+FoTxMnLXWd+79E0J6Rwpdg1BcmZgppjfyHJtY0DWuta7qm5qfTKWvdqesaWmuUZclJ3Z9//snpdp7nZ85txpWT//SzmWlu55o5F8dxGJBSiqmbgFIKQ4tFaQzNQ2uN+XxOyeiJ0LbbLXzfx9PTE2cDBIScuyt9dE0xo08zZtA0zbdPM1JK1pAQAlJKjkMmsKenJ9zd3eH333+HI6XEw8MD3rx5g7/++gsvLy8YjUZc6R2PRzat11RuAuxqpQvGDAUmQIoVBIyeJ6WEbdtwXRdN08BxnLP3+d6psn379i1sAKyRIAjw/v17SClRliVXk12NdE2pm4/1mVrf/fdIn0V0ZbfbndiQ8hpKD/744w/EcYwkSRBFUa/Tmwlln1P+vxP/HjEXjlIgCvS2UgphGEJrje12i19//RXL5ZKTTJrUa5rpSh+g17TWp9G+Z5KYwd28930fSik4tm0jz3PWzmKx4NyHnJL+qc93zPEaMNM/yH9MljODKl2bvQKzmOv2EYBTNRsEwcnMZrMZAHDXIwxDxHHMvTLzZd2J9wE072lifSTQZTfz2mQ8c3SfYQ77w4cPUErBtm1MJhOusff7PZvft0Z31bv35mf3930pkmnS3fd8bT72/f098zoFzjRNuQHXnWB3tYj7qcgys2IKiKaNA3jVB/pM1Bzm//SZuU2Z8nA4hGVZ2Gw2nGpTJDYrwm4K360cu/ddTZirDIDr/654ngfXdXvj02vaccgZpZQYj8eo6xrr9RpVVSGKIs7bKD2noEVpR9M2Zw/smgJVjq9lAN2mYNfZu77U/fsZmKqqcH19jY8fP8K2bVxeXnIznPphpBETDJmBEJp9jibeXf1vgemK+Xt6p/l+8/rMzJIkQZ7nePfuHTzP4zxsNpuhrutelumaVN9LuibZ/R3J10zMbD/1Pc8MHQDgtG3LPWLq8tu2jaIoMJlMsN/vAZyzDiV5SilYUsKCggUF29LAv2LZpw6jsL80MzN+OMKCsHEmjrDgOjY8VwC6RRIPUNc1PDdCHIU4HA4IAw9xNEJd19zrc2zbRlVVGI/HyLIMx+MR19fXsG0bj4+PZy2grlD2IKXkzLYb+c0tjb6O5mvfmY11Kg2on313d4c0TbHb7TCZTKCUwsXFBZzBYIAgCM62KqhPdnNzw/sh3S6k6SNmy5QIhZjH7BP3TbzPFM3rtm2R5znu7u54M6ooCg4l4/EYi8UC6/UaTlEU3FFsmgbj8RhCCHz8+JGrvb4VJM1QWtIVqudd1/2qZqiTSZ90TX5jaobaYLQNcnd3h+fnZ9ze3p7Am1E2z3N4nofFYsFNQZqM2Wgwm3i0CFQ0dZNJSon6FqWvPUtZMPWahRCYzWZQSuFwOODq6gpRFKGqKr53XffUqnJdF6PRCPv9Hp7nIQxDTKdTzOdz1HXNWwpMf8bKmhUfmUy3FOgGzj4wxFwmGGo1UTxr2xZv3rxBFEVYr9cYjUZIkuTU3Pi3aHOapsFqtcIvv/yCh4cHFEWB4/GI29tbaK2xWq3YD0ytEDAa5Cd9YL7mMyYNk7/QDprneUiSBLZt43g8YjAYQEqJOI4xmUyQZRmqqkKSJNjtdnC01oiiCIvFAr7vo2kaJEmC1WrFW319/kCfnucxKCp3+3oAr4Ex41JfrMrzHPf39xgMBsyONzc3eH5+xk8//QQAvBfEuwCUbJLt7/d7CCGw3++xXC5xeXmJzWbDO8uUMZhNdaJmYrKuz3TZ0KRfsntKcsuyRJIkvPustWbHp0ZlkiTn1O+6rqYXEiVmWYb9fs9sQzFHSonBYID1eo3D4cBNCLP11I0zZubd12qSUvKWIRFMmqa4ubnhzSRq11Jco6S4OywAWggBSmvMlVVKYbVaIQxDbLdbnuxut2Pa/Pz5c2+bqVuN9tG7bdsc/Jqmwbt37xggVb1v375FFEVcTcZxDMuyEMcxqEo+A0Pb44PBgNVmmloQBFgul0zf1P3MsgxJkkAp9YVWzHuTCYn1uqwWBAGCIODgO5lMkKYpiqJAmqacxdOi9JUBjuM4qKoKQgg+kBCGITzPw3g85r6ZUgpXV1c8Ga1P2w2bzaa3Z/ZapdhNW+q65i2+x8dHpGnKu2R0rITiEA2tNS4uLnj/iJ+fpqmm/XTzPIq5LU2r8Pfff+P29paj7ufPn2FZFieffZ0YcwX76hc6X0AZ8nQ65bM4o9Hoi15AHMe8l9rrM9R3qqoKw+GQ8x5zErTaQpzOBDw8PHBfresztAAU7L4Gpm1bNi/KBeu6xo8//ojNZoM0TSGEwHA45B0IABxbzsBEUaSLojg7uWS+mHIi+o6OllxcXCDLMqZ0YrPu6O4298Wqm5sbfPr0CT/88AOqquKTTjc3N9jv97yjDID3jABw/nemmS9mYAwCSXufANi/qE9A13mew7ZtlGXJhV63cuyWvJZlIUkS9g+yEvLLbtPiW+Orh+dIXNfVnufpOI41AP3zzz9rnGidD8qtVitN4+XlRZdlqbMs09vtVud5rne7nd7v97ooCn04HHRZllprrZum0VprPkRHz/4/5Os/EEJoIcT5iTvjBB6Bs06HI7SUkkFlWaarqtJVVem6rrWUUjdNc3YikJ7jeR6/z1zA/wXMfwBvwDmgXx7fyAAAAABJRU5ErkJggg=="
             mask="url(#mask4094)"
             id="image4098" />
        </g>
        <path
           d="m 7271,3004.5 c 0,42.2498 -34.25,76.5 -76.5,76.5 -42.25,0 -76.5,-34.2502 -76.5,-76.5 0,-42.2498 34.25,-76.5 76.5,-76.5 42.25,0 76.5,34.2502 76.5,76.5"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4100" />
        <text
           xml:space="preserve"
           transform="matrix(0.75,0,0,-1,7163,2955)"
           style="font-variant:normal;font-weight:normal;font-size:117.875px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text4104"><tspan
             x="0"
             y="0"
             id="tspan4102">V</tspan></text>
      </g>
    </g>
    <g
       id="g4106">
      <g
         id="g4108"
         clip-path="url(#clipPath4112)" />
    </g>
    <g
       id="g4114">
      <g
         id="g4116"
         clip-path="url(#clipPath4120)">
        <g
           id="g4122"
           transform="matrix(153,0,0,153,7024,3108)">
          <image
             width="1"
             height="1"
             style="image-rendering:optimizeSpeed"
             preserveAspectRatio="none"
             transform="matrix(1,0,0,-1,0,1)"
             xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAADMAAAAzCAYAAAA6oTAqAAAABHNCSVQICAgIfAhkiAAADOlJREFUaIGdWllz2zYXPQDBnVopL8qodt3JSx/6//9IO+mD63HcOJIta6EW7iS+B+XCECI76YeZO6JlisTBuRvuBQDI98T3fck5V9f0fRAE6loIIYuikG3bSimlrKpKSillWZaybVvZNI0Sukcf+vs455IxJgFIxpgUQkgAst/vq3fR/01h3y7eHbZto6oqAIAQAk3TQEoJy7JQ1zUeHh5wdXWF3W4H27YBAK7roqoqlGV59CzG2JG4ros0TREEAcIwRJqmAADO+dF99H7LstA0DYIgQFmWqOv69dk/AiOEgOM4SNMUnuehaRq0bYskSRCGobovSRJIKeG6Lvb7PYqiQNM0R/cQGH2ilmXBcRzYto3tdotOpwPP81AUhZo4jfF4jOl0Cs/zkOf5d3P9IRjOOdq2BQCUZYmiKBBFEXa7HaSUuL+/x83NDV5eXhBFERhj2O12YIzB8zyUZQkpJRhjJ8GUZYk4jpEkCQaDATzPQ1VVsG376Bk0h7eA/BQY+rGUEsvlEsPhENvtFnmeg3OOKIqQJAmKokCapmqitm2jrmsURXHEignGcRx0u12lXq7rIgxD1HWNIAjUvaS2bdui1+thu90qgD8NBgDSNIVt27AsCw8PDxgOh8jzHEVRoCxLfPnyBZPJBJvNBkIIMMYgpcR2u4XjOEdACIzJzng8BgDUdY0oihCGIZbLJVzXRa/XU8zSGI1GeHl5+W9gqqqCEAJZlmE6nSKOY2RZhuVyCSGEAtvr9ZAkCdq2RdM0sG0bnHPs9/vvVEwH4/s+wjDEfD6H7/s4Pz/H8/Mzbm5ucHB0B+0gtvv9PubzOQB8Z1M/BCOlxGq1QhRFyPMci8UCeZ6r1U+SBEEQYLFYKHUoigJFUYBzDsuyjpgxwQAHb+m6LpqmQRRF6Pf7mM1muLq6Uk6kaRr4vq9sWAhx5MkAgFmWJUnvyQVzztE0Deq6hpQSRVEgz3NUVaWkLEtUVYWiKFDXNeq6VjospVRSVZVaYQBHYDjncBwHnHMIIWDbtvKerutCCIHz83Os12uMRiNUVYX9fo84jiGEUG6fHJJihr7wPA9ZliHLMrRti7IsUZalspG6rhUI+h+BofhD0rbtcRzQmLEsSzFpWRaEEEoIDIGrqgqj0Qi+78P3fdR1reKZ7m0FAPi+r1AKIbDdbsEYU95IB0Os0DUBqapKxSACQvZjgrEsC5ZlqYnoYGzbVs9omgZxHCu1nk6n6PV6GA6HqKoKnucpb9rpdCDCMMR+vwcAxHGMT58+qXixWq3URE0hVgAolWyaRgEiIWb0IEnM6WD0haD7pZR4enpCHMfY7/fgnKPf7yNJEnS7XTDGkCQJACDLMghKExzHwXQ6hW3beHl5ge/7mM1mcBxHGfQpZmjCpG46I6aa6awQM3RNcUkH1TQNqqpCHMcoyxLdbhebzQaMMWXDZFtpmkKUZQnGGIqiwHw+x263w/n5OR4fHzEYDLBer5Uq6UIsEAhSOZMZU81MMLZtqwyBVJuY4pzj8vIS0+kUUkrYtq1s+urqCk9PTyjL8jWW2bYt67rGdDpFp9NBEAT4999/1cqbNvOWA9BtRhfdk5kOgLwYMUPiui48z4Nt20jTFNfX14iiSKU1v//+O9brNfr9Pnq93muwFkJIMjCK5o7jYL1eI01TpUJ5nh9NXHcApA7kynUgnPN3XTOx9RaYMAxVIur7PobDIdI0xWg0Unmcyj6I1tVqBcYYer2ecrFRFKmciYyc7IBYqOoWdd2gqhrUdaPc5KveVyo4HgDIIxGWBc4ZAA4pGdoWaBqJtgWkZKjrFpYl4boCjFlI0xy+H6r7KMO2bRvCcRysVisMBgPUdY3b21u4rotut4vVaqVUiUT3aAdQrbIfXc3IY5HNmNGfRGqqSL8lthhjEEKAc46qqo5Uk753XVvto8Rms4Hruvj69SviOIbnedhsNmjbVnkOc4K6DRBjBM60GZrcKRXjnEN8S3c450eqSJOlT3I8tCGk6zzPEUURHMeBcF0Xy+USxFCWZej1euCcoyxL7Ha7N2MIeSsS05uR/ehxRjd+xhisb7FGv9/8PPVOunYcB/P5/JD41nUNzjmGwyFmsxmapsFsNkOSJMp2yOBJSN1IzXRQ+gtPgaFB7phcMP2GvntroUzRE1JBuc/9/T3qulZJ3H6/x2Qywf39/VG+pedd5Ax0RvT8jO7RbUbfUFFcMYGSjZB6maqlXwdBAOCwHeCbzQZnZ2eYTCYQQmA+n6sc6fHx8buNlDnMYGqqwY9EZ9R0JPrCEJvmda/Xw93dHQBAdLtdJEmCNE0xGAxQliWyLIOUEt1uFy8vL0dU67naKVvSWaFPWgSTlR8NPWMwgy19TqdT/PbbbyjLEkJKCcdxUNf1kfeifIdWQZ+07nFs+9itmtsAEp1ZeodeD6D30DPIlqmGYGbUNAffP5SnXNcFxxtDf4FpA6e8yinXrWfA9KkzQjbzlqc89W7TKejjCIz+Uv3lppgPfw+Q+UwT1Kn7zXRHZ09fKP1334E5BUTXVV13dWDmQ/Vn6Kt7aiL6xM1NGom+C9VjlAlQmBMxGTn1nb6qZkQ3V49ih/ni97ICc5tgLuBbbIn3gJCh6itpMkeVRz2/IoP/mQzABGcuxnvjXTCnmKAVIuqpJkYT5u2rOlH0NrcB74HR1cdUY52NU6xRGetNZkxQQoiTrhn4Fqnrw98EAjiOJ3rd7NReRrcHE5gp9D/9Xn3wPM/h+76aAOU5bdsiCIKTDz1aXbRgaMGZBGcSFgeExZQ4tqXEFlyJsBhswcE5cGi3tEoYk+Ac4Bxo2xph6KNtaziOQKcToigy1HUJxxFqnkIIiCAIsFwu0e12sd/v8eeffyIMQ1xcXODTp0/fUW1+EnNUddFV7lQuZjJD3kr3Wron8zxP7WCpmjqZTDAYDLDZbDAej/H09ITLy0sIxhiyLFNpyh9//IG///4bt7e3iOMY6/X6JCOWZalMAXjNgs10nrzZ/wuGin7j8Riu66qORJqmSoMuLy9fbcayLHiehzRN8ddff2EymagUhyqHp6I02YfOhglGd9enwLynxmQf9Nwsy47qBWdnZ6oG8PXrVwjf9+E4jspAh8Mh7u7uEAQBVqvVIef5VpQwXSWl4yYY3ZsRGDNGvMcMFTAoFzs/P4eUElmW4fz8HEEQIM9zbDYbdLtdfPny5QA8yzK18owx7Pd7RFGETqeD7XarVupU2qHvy3Ub0bNmvQZwCozneQoAMUHVGao3k0rf3Nyo9ken01FVTSEOjkBQX+X6+hp3d3eqgvjw8ICzszMkSfImM6dyKFPN9C3AKTWjiqTOjOu6R0JdudFohPV6Dc45er2e6ulkWXZ4TpIk8DwPj4+PCIIAdV0jz3NVMSRvRS/Ss1Z9mBnAW0nnqQV4T8qyxPX1NbIsU39/+PAB8/kcHz9+VECKoji0NMjISG3qusZut4NlWdjv93h8fMTl5SXW6zUWiwUuLi4wnU7RNA2yLDvq15BjICB64dzcYDF26GmGYahUpd/vq+52t9uFEEJtjakgSPdGUXTcMrFtW+o9dsuysF6vVcc4CAI0TYPn52dVfCB/T6tilpresplTK19VFfr9vrJbAjQej1EUBaQ8tON934eUEr7vo9PpnMzlGABpWRY6nY6ql9HKtm2L+XwO27aRZRkYO1Tft9stPM+DZVmYzWbfNZv0fc6p3EwXCn51XeP6+loB7PV6mM1mmEwmqgVJ/U/GGMIwBOcc2+32GAzpHJ16AKBUDTi0s5fLJWzbxmKxgOM42Gw2eH5+RhRFqkqjs6K3BXWHQbFFTzrJq9GhCcuyEMexapEPBgMURaGA6Fm6PoQQQp2GoD0/xR4qcFC8GAwGyPNc6exwOFT1NbNrRt+Zmbi5N8nzHKPRCEEQYDqdYjAY4OLiQnWzfd9X3k53NnEcY7FYHKtZv9+X6/VaMUAFBL2jRqvwzz//II5jLJdL/Prrr/j8+bPSdZ0Zs2amgzFTe9d1VfDknOPs7EzZLVVW9b1PGIYnz+QoNXMcB4wdGk7dbhdVVYGCKQ1aZZro09MTXNc92aClBdA3Z2+BIaNumgbj8VgV63/55RfV7uOco9vtKs8JQHXRjsCEYSj3+/3RySX9xY7jqLMqdAJpuVxiNBopQHodzRxm5+wUoA8fPuDz58+4urpCURTwPA/b7Rbj8Rj7/V4dmAAO7Uq9mfyfTjURSP0hZF+O4ygWPc/DbrcD51wdTynL8uShBr0mMBgMVLeYnAFtxU+p0nvjp87OEChiarfb4ePHj7i9vQXweiRlsVggjmMAwGq1UieSzLqCLnRWhvIvWrT/F9C7JwEty5KWZR2fuNNO4umnA6U8nAJ8eXmRUkq5Wq1kURSyKApZlqWsqkrWdX10IpB+6zjOd6cM6RTgz8r/AGeNavoYTAkeAAAAAElFTkSuQmCC"
             mask="url(#mask4124)"
             id="image4128" />
        </g>
        <path
           d="m 7177,3184.5 c 0,42.2498 -34.25,76.5 -76.5,76.5 -42.25,0 -76.5,-34.2502 -76.5,-76.5 0,-42.2498 34.25,-76.5 76.5,-76.5 42.25,0 76.5,34.2502 76.5,76.5"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4130" />
        <text
           xml:space="preserve"
           transform="matrix(0.75,0,0,-1,7068,3135)"
           style="font-variant:normal;font-weight:normal;font-size:117.875px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text4134"><tspan
             x="0"
             y="0"
             id="tspan4132">V</tspan></text>
        <path
           d="m 2402,18933 209,-397"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4136" />
        <path
           d="m 2786,18204 174,-332"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4138" />
        <path
           d="m 3135,17540 174,-332"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4140" />
        <path
           d="m 3483,16876 872,-1660"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4142" />
        <path
           d="m 4530,14884 174,-332"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4144" />
        <path
           d="m 4879,14220 174,-332"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4146" />
        <path
           d="m 5227,13556 872,-1660"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4148" />
        <path
           d="m 6274,11564 174,-332"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4150" />
        <path
           d="m 6623,10900 174,-332"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4152" />
        <path
           d="M 6971,10236 7843,8576"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4154" />
        <path
           d="m 8018,8244 174,-332"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4156" />
        <path
           d="m 8367,7580 174,-332"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4158" />
        <path
           d="M 8715,6916 9587,5256"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4160" />
        <path
           d="m 9762,4924 174,-332"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4162" />
        <path
           d="m 10111,4260 174,-332"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4164" />
        <path
           d="m 10459,3596 951,-1809"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4166" />
        <path
           d="m 11659,1787 469,246 75,-145"
           style="fill:none;stroke:#00dd00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4168" />
        <path
           d="m 2064,18933 81,-154"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4170" />
        <path
           d="m 2319,18447 175,-332"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4172" />
        <path
           d="m 2668,17783 872,-1660"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4174" />
        <path
           d="m 3714,15791 175,-332"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4176" />
        <path
           d="m 4063,15127 175,-332"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4178" />
        <path
           d="m 4412,14463 872,-1660"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4180" />
        <path
           d="m 5458,12471 175,-332"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4182" />
        <path
           d="m 5807,11807 175,-332"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4184" />
        <path
           d="M 6156,11143 7028,9483"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4186" />
        <path
           d="m 7202,9151 175,-332"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4188" />
        <path
           d="m 7551,8487 175,-332"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4190" />
        <path
           d="M 7900,7823 8772,6163"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4192" />
        <path
           d="m 8946,5831 175,-332"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4194" />
        <path
           d="m 9295,5167 175,-332"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4196" />
        <path
           d="m 9644,4503 872,-1660"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4198" />
        <path
           d="m 10690,2511 175,-332"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4200" />
        <path
           d="m 11039,1847 32,-60"
           style="fill:none;stroke:#ff3f00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4202" />
        <path
           d="m 4556,1787 117,30"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4204" />
        <path
           d="m 5035,1914 1443,383"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4206" />
        <path
           d="m 454,4126 1266,336"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4208" />
        <path
           d="m 2083,4558 362,96"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4210" />
        <path
           d="m 2808,4751 362,96"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4212" />
        <path
           d="m 3533,4943 1443,383"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4214" />
        <path
           d="m 454,13277 303,80"
           style="fill:none;stroke:#00bfff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4216" />
        <path
           d="m 11015,4501 -952,-500"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4218" />
        <path
           d="m 9897,3914 -166,-87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4220" />
        <path
           d="m 9565,3739 -166,-87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4222" />
        <path
           d="M 9233,3565 8403,3129"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4224" />
        <path
           d="m 8237,3042 -166,-87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4226" />
        <path
           d="m 7905,2867 -166,-87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4228" />
        <path
           d="M 7573,2693 6621,2193"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4230" />
        <path
           d="M 10714,5076 9761,4576"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4232" />
        <path
           d="m 9596,4488 -166,-87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4234" />
        <path
           d="m 9264,4314 -166,-87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4236" />
        <path
           d="M 8932,4140 8102,3704"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4238" />
        <path
           d="m 7936,3616 -166,-87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4240" />
        <path
           d="m 7604,3442 -166,-87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4242" />
        <path
           d="M 7272,3268 6320,2768"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4244" />
        <path
           d="m 12203,8655 -162,-86"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4246" />
        <path
           d="m 11875,8481 -166,-88"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4248" />
        <path
           d="m 11544,8305 -166,-87"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4250" />
        <path
           d="m 11212,8130 -828,-439"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4252" />
        <path
           d="m 10218,7603 -165,-88"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4254" />
        <path
           d="m 9887,7427 -166,-87"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4256" />
        <path
           d="M 9556,7252 8727,6813"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4258" />
        <path
           d="m 8562,6725 -166,-88"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4260" />
        <path
           d="m 8230,6549 -165,-88"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4262" />
        <path
           d="M 7899,6374 7336,6075 6559,5905"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4264" />
        <path
           d="m 6376,5864 -183,-40"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4266" />
        <path
           d="m 6010,5784 -184,-40"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4268" />
        <path
           d="M 5643,5703 4867,5533"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4270" />
        <path
           d="m 2621,9808 233,122"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4272" />
        <path
           d="m 3020,10017 332,174"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4274" />
        <path
           d="m 3518,10278 332,175"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4276" />
        <path
           d="m 4016,10540 332,174"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4278" />
        <path
           d="m 4514,10802 332,174"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4280" />
        <path
           d="m 5012,11063 332,175"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4282" />
        <path
           d="m 5510,11325 332,174"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4284" />
        <path
           d="m 6008,11586 332,175"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4286" />
        <path
           d="m 6506,11848 332,174"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4288" />
        <path
           d="m 7004,12110 332,174"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4290" />
        <path
           d="m 7502,12371 332,175"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4292" />
        <path
           d="m 8000,12633 332,174"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4294" />
        <path
           d="m 8498,12894 332,175"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4296" />
        <path
           d="m 8996,13156 332,174"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4298" />
        <path
           d="m 9494,13418 332,174"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4300" />
        <path
           d="m 9992,13679 332,175"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4302" />
        <path
           d="m 10490,13941 332,174"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4304" />
        <path
           d="m 10988,14202 332,175"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4306" />
        <path
           d="m 11486,14464 232,122"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4308" />
        <path
           d="m 7205,11754 808,425"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4310" />
        <path
           d="m 8179,12266 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4312" />
        <path
           d="m 8511,12440 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4314" />
        <path
           d="m 8843,12615 830,436"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4316" />
        <path
           d="m 9839,13138 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4318" />
        <path
           d="m 10171,13312 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4320" />
        <path
           d="m 10503,13487 830,436"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4322" />
        <path
           d="m 11499,14010 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4324" />
        <path
           d="m 11831,14184 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4326" />
        <path
           d="m 12163,14359 40,21"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4328" />
        <path
           d="m 6770,12583 807,424"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4330" />
        <path
           d="m 7743,13094 166,88"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4332" />
        <path
           d="m 8075,13269 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4334" />
        <path
           d="m 8407,13443 830,436"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4336" />
        <path
           d="m 9403,13966 166,88"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4338" />
        <path
           d="m 9735,14141 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4340" />
        <path
           d="m 10067,14315 830,436"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4342" />
        <path
           d="m 11063,14838 166,88"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4344" />
        <path
           d="m 11395,15013 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4346" />
        <path
           d="m 11727,15187 476,250"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4348" />
        <path
           d="m 4683,9108 532,279 -279,531 -532,-279 279,-531"
           style="fill:none;stroke:#0000ff;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4350" />
        <path
           d="m 4217.5698,9562.7344 c -89.2593,-44.3096 -135.9944,-144.4727 -112.6064,-241.3418 23.3877,-96.8682 110.6767,-164.6738 210.3203,-163.374"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4352" />
        <path
           d="m 4315.5127,9157.9297 c -52.9902,-96.6709 -27.5772,-217.5401 59.8555,-284.6875 87.4326,-67.1475 210.7666,-60.5137 290.4921,15.625"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4354" />
        <path
           d="m 4664.7812,8889.1445 c 25.8389,-98.0722 119.3614,-162.6289 220.2237,-152.0166 100.8623,10.6133 178.8994,93.2227 183.7593,194.5244"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4356" />
        <path
           d="m 5069.3071,8931.7197 c 68.1529,-55.8115 167.1197,-52.4541 231.333,7.8487 64.2134,60.3027 73.7754,158.8632 22.3511,230.3847"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4358" />
        <path
           d="m 5323.5019,9171.0059 c 128.9273,-17.6993 255.9087,43.58 322.2725,155.5224 66.3643,111.9434 59.1895,252.7549 -18.209,357.3731 -77.3984,104.6181 -209.9507,152.6728 -336.4111,121.9609"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4360" />
        <path
           d="m 5291.0669,9806.3691 c 37.9609,55.4219 42.4062,127.2178 11.5723,186.8995 -30.8345,59.6814 -91.9629,97.5984 -159.1299,98.7074"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4362" />
        <path
           d="m 5143.8945,10091.776 c -44.9751,157.115 -203.1001,253.325 -363.3066,221.05 -160.207,-32.274 -268.7461,-182.205 -249.3789,-344.4783"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4364" />
        <path
           d="m 4531.4204,9967.4492 c -112.2461,77.6438 -265.6362,53.7918 -349.0059,-54.2695 -83.3691,-108.0615 -67.5166,-262.4834 36.0689,-351.3526"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path4366" />
        <path
           d="m 5466,5199 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4368" />
        <path
           d="m 6332,5348 -17,4"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4370" />
        <path
           d="m 5835,5471 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4372" />
        <path
           d="m 5311,5602 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4374" />
        <path
           d="m 4787,5733 -29,7"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4376" />
        <path
           d="m 6728,5614 -43,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4378" />
        <path
           d="m 6204,5744 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4380" />
        <path
           d="m 5680,5875 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4382" />
        <path
           d="m 5156,6005 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4384" />
        <path
           d="m 4632,6136 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4386" />
        <path
           d="m 6573,6017 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4388" />
        <path
           d="m 6049,6147 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4390" />
        <path
           d="m 5526,6278 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4392" />
        <path
           d="m 5002,6409 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4394" />
        <path
           d="m 5895,6551 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4396" />
        <path
           d="m 5371,6681 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4398" />
        <path
           d="m 4847,6812 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4400" />
        <path
           d="m 5740,6954 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4402" />
        <path
           d="m 5216,7085 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4404" />
        <path
           d="m 4692,7215 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4406" />
        <path
           d="m 4168,7346 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4408" />
        <path
           d="m 5585,7357 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4410" />
        <path
           d="m 5061,7488 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4412" />
        <path
           d="m 4537,7619 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4414" />
        <path
           d="m 4013,7749 -37,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4416" />
        <path
           d="m 5949,7631 -38,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4418" />
        <path
           d="m 5430,7761 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4420" />
        <path
           d="m 4906,7891 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4422" />
        <path
           d="m 4382,8022 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4424" />
        <path
           d="m 3858,8153 -33,8"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4426" />
        <path
           d="m 5799,8033 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4428" />
        <path
           d="m 5275,8164 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4430" />
        <path
           d="m 4751,8295 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4432" />
        <path
           d="m 4227,8425 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4434" />
        <path
           d="m 3703,8556 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4436" />
        <path
           d="m 5645,8437 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4438" />
        <path
           d="m 3025,9090 -31,7"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4440" />
        <path
           d="m 5121,8567 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4442" />
        <path
           d="m 4597,8698 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4444" />
        <path
           d="m 4073,8829 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4446" />
        <path
           d="m 3549,8959 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4448" />
        <path
           d="m 5490,8840 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4450" />
        <path
           d="m 2870,9493 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4452" />
        <path
           d="m 4442,9101 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4454" />
        <path
           d="m 3918,9232 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4456" />
        <path
           d="m 3394,9363 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4458" />
        <path
           d="m 2715,9897 -44,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4460" />
        <path
           d="m 4287,9505 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4462" />
        <path
           d="m 3763,9635 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4464" />
        <path
           d="m 3239,9766 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4466" />
        <path
           d="m 4656,9777 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4468" />
        <path
           d="m 4132,9908 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4470" />
        <path
           d="m 3608,10039 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4472" />
        <path
           d="m 3084,10169 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4474" />
        <path
           d="m 2560,10300 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4476" />
        <path
           d="m 4501,10181 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4478" />
        <path
           d="m 3977,10311 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4480" />
        <path
           d="m 3453,10442 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4482" />
        <path
           d="m 2929,10573 -43,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4484" />
        <path
           d="m 2405,10703 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4486" />
        <path
           d="m 4346,10584 -3,1"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4488" />
        <path
           d="m 3823,10715 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4490" />
        <path
           d="m 3299,10845 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4492" />
        <path
           d="m 2775,10976 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4494" />
        <path
           d="m 2251,11107 -44,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4496" />
        <path
           d="m 4192,10987 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4498" />
        <path
           d="m 3668,11118 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4500" />
        <path
           d="m 3144,11249 -44,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4502" />
        <path
           d="m 2620,11379 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4504" />
        <path
           d="m 2096,11510 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4506" />
        <path
           d="m 4037,11391 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4508" />
        <path
           d="m 3513,11521 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4510" />
        <path
           d="m 2989,11652 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4512" />
        <path
           d="m 2465,11783 -44,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4514" />
        <path
           d="m 1941,11913 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4516" />
        <path
           d="m 3882,11794 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4518" />
        <path
           d="m 3358,11925 -44,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4520" />
        <path
           d="m 2834,12055 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4522" />
        <path
           d="m 2310,12186 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4524" />
        <path
           d="m 1786,12317 -44,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4526" />
        <path
           d="m 1262,12447 -31,8"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4528" />
        <path
           d="m 3727,12197 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4530" />
        <path
           d="m 3203,12328 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4532" />
        <path
           d="m 2679,12459 -43,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4534" />
        <path
           d="m 2155,12589 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4536" />
        <path
           d="m 1631,12720 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4538" />
        <path
           d="m 1107,12850 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4540" />
        <path
           d="m 3048,12731 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4542" />
        <path
           d="m 2524,12862 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4544" />
        <path
           d="m 2000,12992 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4546" />
        <path
           d="m 1476,13123 -43,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4548" />
        <path
           d="m 953,13254 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4550" />
        <path
           d="m 2894,13135 -44,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4552" />
        <path
           d="m 2370,13265 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4554" />
        <path
           d="m 1846,13396 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4556" />
        <path
           d="m 1322,13526 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4558" />
        <path
           d="m 798,13657 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4560" />
        <path
           d="m 2739,13538 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4562" />
        <path
           d="m 2215,13668 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4564" />
        <path
           d="m 1691,13799 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4566" />
        <path
           d="m 1167,13930 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4568" />
        <path
           d="m 2584,13941 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4570" />
        <path
           d="m 2060,14072 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4572" />
        <path
           d="m 1536,14202 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4574" />
        <path
           d="m 1905,14475 -44,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4576" />
        <path
           d="m 1262,12447 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4578" />
        <path
           d="m 1107,12850 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4580" />
        <path
           d="m 953,13254 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4582" />
        <path
           d="m 798,13657 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4584" />
        <path
           d="m 3025,9090 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4586" />
        <path
           d="m 2870,9493 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4588" />
        <path
           d="m 2715,9897 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4590" />
        <path
           d="m 2560,10300 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4592" />
        <path
           d="m 2405,10703 -12,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4594" />
        <path
           d="m 2251,11107 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4596" />
        <path
           d="m 2096,11510 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4598" />
        <path
           d="m 1941,11913 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4600" />
        <path
           d="m 1786,12317 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4602" />
        <path
           d="m 1631,12720 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4604" />
        <path
           d="m 1476,13123 -12,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4606" />
        <path
           d="m 1322,13526 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4608" />
        <path
           d="m 1167,13930 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4610" />
        <path
           d="m 4787,5733 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4612" />
        <path
           d="m 4632,6136 -6,17"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4614" />
        <path
           d="m 3858,8153 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4616" />
        <path
           d="m 3703,8556 -12,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4618" />
        <path
           d="m 3549,8959 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4620" />
        <path
           d="m 3394,9363 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4622" />
        <path
           d="m 3239,9766 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4624" />
        <path
           d="m 3084,10169 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4626" />
        <path
           d="m 2929,10573 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4628" />
        <path
           d="m 2775,10976 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4630" />
        <path
           d="m 2620,11379 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4632" />
        <path
           d="m 2465,11783 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4634" />
        <path
           d="m 2310,12186 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4636" />
        <path
           d="m 2155,12589 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4638" />
        <path
           d="m 2000,12992 -12,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4640" />
        <path
           d="m 1846,13396 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4642" />
        <path
           d="m 1691,13799 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4644" />
        <path
           d="m 1536,14202 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4646" />
        <path
           d="m 4168,7346 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4648" />
        <path
           d="m 4013,7749 -9,24"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4650" />
        <path
           d="m 5466,5199 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4652" />
        <path
           d="m 5311,5602 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4654" />
        <path
           d="m 5156,6005 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4656" />
        <path
           d="m 5002,6409 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4658" />
        <path
           d="m 4847,6812 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4660" />
        <path
           d="m 4692,7215 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4662" />
        <path
           d="m 4537,7619 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4664" />
        <path
           d="m 1905,14475 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4666" />
        <path
           d="m 4382,8022 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4668" />
        <path
           d="m 4227,8425 -12,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4670" />
        <path
           d="m 4073,8829 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4672" />
        <path
           d="m 3918,9232 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4674" />
        <path
           d="m 3763,9635 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4676" />
        <path
           d="m 3608,10039 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4678" />
        <path
           d="m 3453,10442 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4680" />
        <path
           d="m 3299,10845 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4682" />
        <path
           d="m 3144,11249 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4684" />
        <path
           d="m 2989,11652 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4686" />
        <path
           d="m 2834,12055 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4688" />
        <path
           d="m 2679,12459 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4690" />
        <path
           d="m 2524,12862 -12,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4692" />
        <path
           d="m 2370,13265 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4694" />
        <path
           d="m 2215,13668 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4696" />
        <path
           d="m 2060,14072 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4698" />
        <path
           d="m 5835,5471 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4700" />
        <path
           d="m 5680,5875 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4702" />
        <path
           d="m 5526,6278 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4704" />
        <path
           d="m 5371,6681 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4706" />
        <path
           d="m 5216,7085 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4708" />
        <path
           d="m 5061,7488 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4710" />
        <path
           d="m 4906,7891 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4712" />
        <path
           d="m 4751,8295 -12,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4714" />
        <path
           d="m 4597,8698 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4716" />
        <path
           d="m 4442,9101 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4718" />
        <path
           d="m 4287,9505 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4720" />
        <path
           d="m 4132,9908 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4722" />
        <path
           d="m 3977,10311 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4724" />
        <path
           d="m 3823,10715 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4726" />
        <path
           d="m 3668,11118 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4728" />
        <path
           d="m 3513,11521 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4730" />
        <path
           d="m 3358,11925 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4732" />
        <path
           d="m 3203,12328 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4734" />
        <path
           d="m 3048,12731 -12,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4736" />
        <path
           d="m 2894,13135 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4738" />
        <path
           d="m 2739,13538 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4740" />
        <path
           d="m 2584,13941 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4742" />
        <path
           d="m 6355,5353 -9,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4744" />
        <path
           d="m 6204,5744 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4746" />
        <path
           d="m 6049,6147 -12,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4748" />
        <path
           d="m 5895,6551 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4750" />
        <path
           d="m 5740,6954 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4752" />
        <path
           d="m 5585,7357 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4754" />
        <path
           d="m 5430,7761 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4756" />
        <path
           d="m 5275,8164 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4758" />
        <path
           d="m 5121,8567 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4760" />
        <path
           d="m 4192,10987 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4762" />
        <path
           d="m 4037,11391 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4764" />
        <path
           d="m 3882,11794 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4766" />
        <path
           d="m 3727,12197 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4768" />
        <path
           d="m 4656,9777 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4770" />
        <path
           d="m 4501,10181 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4772" />
        <path
           d="m 4346,10584 v 2"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4774" />
        <path
           d="m 6728,5614 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4776" />
        <path
           d="m 6573,6017 -12,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4778" />
        <path
           d="m 5953,7634 -12,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4780" />
        <path
           d="m 5799,8033 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4782" />
        <path
           d="m 5645,8437 -13,33"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4784" />
        <path
           d="m 5490,8840 -13,34"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4786" />
        <path
           d="m 6715,5647 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4788" />
        <path
           d="m 6346,5374 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4790" />
        <path
           d="m 6561,6050 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4792" />
        <path
           d="m 6191,5778 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4794" />
        <path
           d="m 5822,5505 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4796" />
        <path
           d="m 5453,5232 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4798" />
        <path
           d="m 6037,6181 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4800" />
        <path
           d="m 5667,5908 -30,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4802" />
        <path
           d="m 5298,5636 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4804" />
        <path
           d="m 5882,6584 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4806" />
        <path
           d="m 5513,6312 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4808" />
        <path
           d="m 5143,6039 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4810" />
        <path
           d="m 4774,5766 -21,-16"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4812" />
        <path
           d="m 4618,6168 -29,-21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4814" />
        <path
           d="m 5727,6988 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4816" />
        <path
           d="m 5358,6715 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4818" />
        <path
           d="m 4989,6442 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4820" />
        <path
           d="m 5941,7664 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4822" />
        <path
           d="m 5572,7391 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4824" />
        <path
           d="m 5203,7118 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4826" />
        <path
           d="m 4834,6846 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4828" />
        <path
           d="m 5786,8067 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4830" />
        <path
           d="m 5417,7794 -30,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4832" />
        <path
           d="m 5048,7522 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4834" />
        <path
           d="m 4679,7249 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4836" />
        <path
           d="m 5632,8470 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4838" />
        <path
           d="m 5263,8198 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4840" />
        <path
           d="m 4893,7925 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4842" />
        <path
           d="m 4524,7652 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4844" />
        <path
           d="m 4155,7380 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4846" />
        <path
           d="m 5477,8874 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4848" />
        <path
           d="m 5108,8601 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4850" />
        <path
           d="m 4739,8328 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4852" />
        <path
           d="m 4369,8056 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4854" />
        <path
           d="m 4584,8732 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4856" />
        <path
           d="m 4215,8459 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4858" />
        <path
           d="m 3845,8186 -24,-18"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4860" />
        <path
           d="m 4429,9135 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4862" />
        <path
           d="m 4060,8862 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4864" />
        <path
           d="m 3691,8590 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4866" />
        <path
           d="m 4643,9811 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4868" />
        <path
           d="m 4274,9538 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4870" />
        <path
           d="m 3905,9266 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4872" />
        <path
           d="m 3536,8993 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4874" />
        <path
           d="m 4488,10214 -30,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4876" />
        <path
           d="m 4119,9942 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4878" />
        <path
           d="m 3750,9669 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4880" />
        <path
           d="m 3381,9396 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4882" />
        <path
           d="m 3012,9124 -23,-17"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4884" />
        <path
           d="m 3964,10345 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4886" />
        <path
           d="m 3595,10072 -30,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4888" />
        <path
           d="m 3226,9800 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4890" />
        <path
           d="m 2857,9527 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4892" />
        <path
           d="m 4179,11021 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4894" />
        <path
           d="m 3810,10748 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4896" />
        <path
           d="m 3440,10476 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4898" />
        <path
           d="m 3071,10203 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4900" />
        <path
           d="m 2702,9930 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4902" />
        <path
           d="m 4024,11424 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4904" />
        <path
           d="m 3655,11152 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4906" />
        <path
           d="m 3286,10879 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4908" />
        <path
           d="m 2916,10606 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4910" />
        <path
           d="m 2547,10334 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4912" />
        <path
           d="m 3869,11828 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4914" />
        <path
           d="m 3500,11555 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4916" />
        <path
           d="m 3131,11282 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4918" />
        <path
           d="m 2762,11010 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4920" />
        <path
           d="m 2393,10737 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4922" />
        <path
           d="m 3714,12231 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4924" />
        <path
           d="m 3345,11958 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4926" />
        <path
           d="m 2976,11686 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4928" />
        <path
           d="m 2607,11413 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4930" />
        <path
           d="m 2238,11140 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4932" />
        <path
           d="m 3190,12362 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4934" />
        <path
           d="m 2821,12089 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4936" />
        <path
           d="m 2452,11816 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4938" />
        <path
           d="m 2083,11543 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4940" />
        <path
           d="m 3036,12765 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4942" />
        <path
           d="m 2666,12492 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4944" />
        <path
           d="m 2297,12219 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4946" />
        <path
           d="m 1928,11947 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4948" />
        <path
           d="m 2881,13168 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4950" />
        <path
           d="m 2512,12895 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4952" />
        <path
           d="m 2142,12623 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4954" />
        <path
           d="m 1773,12350 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4956" />
        <path
           d="m 2726,13571 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4958" />
        <path
           d="m 2357,13299 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4960" />
        <path
           d="m 1988,13026 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4962" />
        <path
           d="m 1618,12753 -30,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4964" />
        <path
           d="m 1249,12481 -23,-17"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4966" />
        <path
           d="m 2571,13975 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4968" />
        <path
           d="m 2202,13702 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4970" />
        <path
           d="m 1833,13429 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4972" />
        <path
           d="m 1464,13157 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4974" />
        <path
           d="m 1094,12884 -30,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4976" />
        <path
           d="m 2047,14105 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4978" />
        <path
           d="m 1678,13833 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4980" />
        <path
           d="m 1309,13560 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4982" />
        <path
           d="m 940,13287 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4984" />
        <path
           d="m 1892,14509 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4986" />
        <path
           d="m 1523,14236 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4988" />
        <path
           d="m 1154,13963 -31,-22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4990" />
        <path
           d="m 785,13691 -31,-23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4992" />
        <path
           d="m 5923,5292 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4994" />
        <path
           d="m 5152,5540 -64,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4996" />
        <path
           d="m 6503,5663 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path4998" />
        <path
           d="m 5732,5911 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5000" />
        <path
           d="m 4961,6159 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5002" />
        <path
           d="m 5541,6530 -65,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5004" />
        <path
           d="m 4769,6778 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5006" />
        <path
           d="m 5349,7149 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5008" />
        <path
           d="m 4578,7397 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5010" />
        <path
           d="m 3807,7645 -60,19"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5012" />
        <path
           d="m 5158,7768 -65,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5014" />
        <path
           d="m 4386,8016 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5016" />
        <path
           d="m 5737,8140 -64,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5018" />
        <path
           d="m 4966,8387 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5020" />
        <path
           d="m 4195,8635 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5022" />
        <path
           d="m 3424,8883 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5024" />
        <path
           d="m 5544,8759 -62,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5026" />
        <path
           d="m 4775,9007 -65,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5028" />
        <path
           d="m 4004,9254 -65,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5030" />
        <path
           d="m 3812,9873 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5032" />
        <path
           d="m 3041,10121 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5034" />
        <path
           d="m 4392,10245 -64,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5036" />
        <path
           d="m 3621,10493 -65,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5038" />
        <path
           d="m 2849,10740 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5040" />
        <path
           d="m 2078,10988 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5042" />
        <path
           d="m 4200,10864 -64,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5044" />
        <path
           d="m 3429,11112 -64,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5046" />
        <path
           d="m 2658,11359 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5048" />
        <path
           d="m 1887,11607 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5050" />
        <path
           d="m 4009,11483 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5052" />
        <path
           d="m 3238,11731 -64,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5054" />
        <path
           d="m 2467,11979 -65,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5056" />
        <path
           d="m 1695,12226 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5058" />
        <path
           d="m 3782,12113 -29,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5060" />
        <path
           d="m 3046,12350 -64,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5062" />
        <path
           d="m 2275,12598 -64,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5064" />
        <path
           d="m 1504,12845 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5066" />
        <path
           d="m 2855,12969 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5068" />
        <path
           d="m 2084,13217 -65,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5070" />
        <path
           d="m 1313,13465 -65,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5072" />
        <path
           d="m 2663,13588 -64,21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5074" />
        <path
           d="m 1892,13836 -64,20"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5076" />
        <path
           d="m 1121,14084 -54,17"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5078" />
        <path
           d="m 6488,5715 -49,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5080" />
        <path
           d="m 5908,5343 -48,-30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5082" />
        <path
           d="m 5716,5963 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5084" />
        <path
           d="m 5137,5591 -49,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5086" />
        <path
           d="m 5525,6582 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5088" />
        <path
           d="m 4945,6210 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5090" />
        <path
           d="m 5333,7201 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5092" />
        <path
           d="m 4754,6829 -49,-30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5094" />
        <path
           d="m 5722,8191 -49,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5096" />
        <path
           d="m 5142,7820 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5098" />
        <path
           d="m 4562,7449 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5100" />
        <path
           d="m 5521,8804 -39,-25"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5102" />
        <path
           d="m 3791,7696 -45,-29"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5104" />
        <path
           d="m 4951,8439 -49,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5106" />
        <path
           d="m 4371,8068 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5108" />
        <path
           d="m 4759,9058 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5110" />
        <path
           d="m 4179,8687 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5112" />
        <path
           d="m 3988,9306 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5114" />
        <path
           d="m 3408,8935 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5116" />
        <path
           d="m 4376,10296 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5118" />
        <path
           d="m 3796,9925 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5120" />
        <path
           d="m 4185,10915 -49,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5122" />
        <path
           d="m 3605,10544 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5124" />
        <path
           d="m 3025,10173 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5126" />
        <path
           d="m 3993,11534 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5128" />
        <path
           d="m 3414,11163 -49,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5130" />
        <path
           d="m 2834,10792 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5132" />
        <path
           d="m 3771,12134 -17,-11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5134" />
        <path
           d="m 3222,11782 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5136" />
        <path
           d="m 2642,11411 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5138" />
        <path
           d="m 2063,11040 -49,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5140" />
        <path
           d="m 3031,12401 -49,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5142" />
        <path
           d="m 2451,12030 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5144" />
        <path
           d="m 1871,11659 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5146" />
        <path
           d="m 2839,13020 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5148" />
        <path
           d="m 2259,12649 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5150" />
        <path
           d="m 1680,12278 -49,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5152" />
        <path
           d="m 2648,13639 -49,-30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5154" />
        <path
           d="m 2068,13268 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5156" />
        <path
           d="m 1488,12897 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5158" />
        <path
           d="m 1877,13887 -49,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5160" />
        <path
           d="m 1297,13516 -48,-31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5162" />
        <path
           d="m 2079,10988 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5164" />
        <path
           d="m 1887,11607 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5166" />
        <path
           d="m 1696,12226 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5168" />
        <path
           d="m 1504,12845 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5170" />
        <path
           d="m 1313,13464 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5172" />
        <path
           d="m 1121,14084 -12,39"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5174" />
        <path
           d="m 3807,7645 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5176" />
        <path
           d="m 3041,10121 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5178" />
        <path
           d="m 2850,10740 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5180" />
        <path
           d="m 2658,11359 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5182" />
        <path
           d="m 2467,11978 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5184" />
        <path
           d="m 2275,12598 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5186" />
        <path
           d="m 2084,13217 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5188" />
        <path
           d="m 1893,13836 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5190" />
        <path
           d="m 3424,8883 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5192" />
        <path
           d="m 4387,8016 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5194" />
        <path
           d="m 4195,8635 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5196" />
        <path
           d="m 4004,9254 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5198" />
        <path
           d="m 3812,9873 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5200" />
        <path
           d="m 3621,10492 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5202" />
        <path
           d="m 3430,11112 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5204" />
        <path
           d="m 3238,11731 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5206" />
        <path
           d="m 3047,12350 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5208" />
        <path
           d="m 2855,12969 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5210" />
        <path
           d="m 2664,13588 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5212" />
        <path
           d="m 5153,5540 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5214" />
        <path
           d="m 4961,6159 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5216" />
        <path
           d="m 4770,6778 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5218" />
        <path
           d="m 4578,7397 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5220" />
        <path
           d="m 5924,5292 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5222" />
        <path
           d="m 5732,5911 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5224" />
        <path
           d="m 5541,6530 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5226" />
        <path
           d="m 5349,7149 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5228" />
        <path
           d="m 5158,7768 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5230" />
        <path
           d="m 4967,8387 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5232" />
        <path
           d="m 4775,9006 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5234" />
        <path
           d="m 4201,10864 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5236" />
        <path
           d="m 4009,11483 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5238" />
        <path
           d="m 4392,10245 -16,51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5240" />
        <path
           d="m 6504,5663 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5242" />
        <path
           d="m 5738,8139 -16,52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5244" />
        <path
           d="m 5278,5479 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5246" />
        <path
           d="m 4883,5847 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5248" />
        <path
           d="m 5733,5538 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5250" />
        <path
           d="m 5338,5907 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5252" />
        <path
           d="m 4943,6275 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5254" />
        <path
           d="m 4153,7012 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5256" />
        <path
           d="m 4516,6673 -1,1"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5258" />
        <path
           d="m 6188,5598 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5260" />
        <path
           d="m 5793,5966 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5262" />
        <path
           d="m 5398,6334 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5264" />
        <path
           d="m 5003,6703 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5266" />
        <path
           d="m 4608,7071 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5268" />
        <path
           d="m 4213,7439 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5270" />
        <path
           d="m 6643,5657 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5272" />
        <path
           d="m 6248,6026 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5274" />
        <path
           d="m 5853,6394 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5276" />
        <path
           d="m 5458,6762 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5278" />
        <path
           d="m 5063,7131 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5280" />
        <path
           d="m 4668,7499 -32,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5282" />
        <path
           d="m 4273,7867 -32,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5284" />
        <path
           d="m 3879,8235 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5286" />
        <path
           d="m 3089,8972 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5288" />
        <path
           d="m 3484,8604 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5290" />
        <path
           d="m 7098,5717 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5292" />
        <path
           d="m 6703,6085 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5294" />
        <path
           d="m 2754,9768 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5296" />
        <path
           d="m 5913,6822 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5298" />
        <path
           d="m 5518,7190 -32,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5300" />
        <path
           d="m 5123,7558 -32,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5302" />
        <path
           d="m 4729,7927 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5304" />
        <path
           d="m 4334,8295 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5306" />
        <path
           d="m 3939,8663 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5308" />
        <path
           d="m 3544,9032 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5310" />
        <path
           d="m 6368,6881 -32,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5312" />
        <path
           d="m 5579,7618 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5314" />
        <path
           d="m 5184,7986 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5316" />
        <path
           d="m 4789,8354 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5318" />
        <path
           d="m 4394,8723 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5320" />
        <path
           d="m 3999,9091 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5322" />
        <path
           d="m 3604,9459 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5324" />
        <path
           d="m 3209,9828 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5326" />
        <path
           d="m 2814,10196 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5328" />
        <path
           d="m 2419,10564 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5330" />
        <path
           d="m 6034,7677 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5332" />
        <path
           d="m 5639,8046 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5334" />
        <path
           d="m 4849,8782 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5336" />
        <path
           d="m 4454,9151 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5338" />
        <path
           d="m 4059,9519 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5340" />
        <path
           d="m 3664,9887 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5342" />
        <path
           d="m 3269,10255 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5344" />
        <path
           d="m 2874,10624 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5346" />
        <path
           d="m 2479,10992 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5348" />
        <path
           d="m 2084,11360 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5350" />
        <path
           d="m 1689,11729 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5352" />
        <path
           d="m 5690,8482 -24,22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5354" />
        <path
           d="m 4119,9947 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5356" />
        <path
           d="m 3724,10315 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5358" />
        <path
           d="m 3329,10683 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5360" />
        <path
           d="m 2934,11052 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5362" />
        <path
           d="m 2539,11420 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5364" />
        <path
           d="m 2144,11788 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5366" />
        <path
           d="m 1749,12156 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5368" />
        <path
           d="m 1354,12525 -32,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5370" />
        <path
           d="m 4909,9210 -11,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5372" />
        <path
           d="m 4574,10006 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5374" />
        <path
           d="m 4179,10374 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5376" />
        <path
           d="m 3784,10743 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5378" />
        <path
           d="m 3389,11111 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5380" />
        <path
           d="m 2994,11479 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5382" />
        <path
           d="m 2599,11848 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5384" />
        <path
           d="m 2204,12216 -32,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5386" />
        <path
           d="m 1810,12584 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5388" />
        <path
           d="m 1415,12953 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5390" />
        <path
           d="m 1020,13321 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5392" />
        <path
           d="m 625,13689 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5394" />
        <path
           d="m 4634,10434 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5396" />
        <path
           d="m 4239,10802 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5398" />
        <path
           d="m 3844,11171 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5400" />
        <path
           d="m 3449,11539 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5402" />
        <path
           d="m 3054,11907 -32,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5404" />
        <path
           d="m 2660,12275 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5406" />
        <path
           d="m 2265,12644 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5408" />
        <path
           d="m 1870,13012 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5410" />
        <path
           d="m 1475,13380 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5412" />
        <path
           d="m 1080,13749 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5414" />
        <path
           d="m 3904,11598 -32,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5416" />
        <path
           d="m 3510,11967 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5418" />
        <path
           d="m 3115,12335 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5420" />
        <path
           d="m 2720,12703 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5422" />
        <path
           d="m 2325,13072 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5424" />
        <path
           d="m 1930,13440 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5426" />
        <path
           d="m 1535,13808 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5428" />
        <path
           d="m 3570,12395 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5430" />
        <path
           d="m 3175,12763 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5432" />
        <path
           d="m 2780,13131 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5434" />
        <path
           d="m 2385,13499 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5436" />
        <path
           d="m 1990,13868 -33,30"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5438" />
        <path
           d="m 1595,14236 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5440" />
        <path
           d="m 2840,13559 -33,31"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5442" />
        <path
           d="m 2445,13927 -23,22"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5444" />
        <path
           d="m 625,13689 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5446" />
        <path
           d="m 1020,13321 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5448" />
        <path
           d="m 1080,13749 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5450" />
        <path
           d="m 1354,12525 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5452" />
        <path
           d="m 1415,12953 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5454" />
        <path
           d="m 1475,13380 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5456" />
        <path
           d="m 1535,13808 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5458" />
        <path
           d="m 1595,14236 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5460" />
        <path
           d="m 1689,11729 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5462" />
        <path
           d="m 1749,12156 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5464" />
        <path
           d="m 1810,12584 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5466" />
        <path
           d="m 1870,13012 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5468" />
        <path
           d="m 1930,13440 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5470" />
        <path
           d="m 1990,13868 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5472" />
        <path
           d="m 2025,10942 4,26"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5474" />
        <path
           d="m 2084,11360 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5476" />
        <path
           d="m 2144,11788 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5478" />
        <path
           d="m 2204,12216 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5480" />
        <path
           d="m 2265,12644 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5482" />
        <path
           d="m 2325,13072 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5484" />
        <path
           d="m 2385,13499 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5486" />
        <path
           d="m 2445,13927 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5488" />
        <path
           d="m 2419,10564 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5490" />
        <path
           d="m 2479,10992 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5492" />
        <path
           d="m 2539,11420 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5494" />
        <path
           d="m 2599,11848 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5496" />
        <path
           d="m 2660,12275 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5498" />
        <path
           d="m 2720,12703 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5500" />
        <path
           d="m 2780,13131 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5502" />
        <path
           d="m 2840,13559 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5504" />
        <path
           d="m 2754,9768 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5506" />
        <path
           d="m 2814,10196 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5508" />
        <path
           d="m 2874,10624 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5510" />
        <path
           d="m 2934,11052 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5512" />
        <path
           d="m 2994,11479 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5514" />
        <path
           d="m 3054,11907 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5516" />
        <path
           d="m 3115,12335 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5518" />
        <path
           d="m 3175,12763 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5520" />
        <path
           d="m 3089,8972 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5522" />
        <path
           d="m 3209,9828 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5524" />
        <path
           d="m 3269,10255 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5526" />
        <path
           d="m 3329,10683 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5528" />
        <path
           d="m 3389,11111 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5530" />
        <path
           d="m 3449,11539 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5532" />
        <path
           d="m 3510,11967 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5534" />
        <path
           d="m 3570,12395 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5536" />
        <path
           d="m 3484,8604 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5538" />
        <path
           d="m 3544,9032 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5540" />
        <path
           d="m 3604,9459 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5542" />
        <path
           d="m 3664,9887 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5544" />
        <path
           d="m 3724,10315 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5546" />
        <path
           d="m 3784,10743 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5548" />
        <path
           d="m 3844,11171 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5550" />
        <path
           d="m 3904,11598 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5552" />
        <path
           d="m 4239,10802 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5554" />
        <path
           d="m 3879,8235 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5556" />
        <path
           d="m 3939,8663 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5558" />
        <path
           d="m 3999,9091 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5560" />
        <path
           d="m 4059,9519 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5562" />
        <path
           d="m 4119,9947 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5564" />
        <path
           d="m 4179,10374 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5566" />
        <path
           d="m 4153,7012 5,32"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5568" />
        <path
           d="m 4574,10006 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5570" />
        <path
           d="m 4634,10434 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5572" />
        <path
           d="m 4213,7439 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5574" />
        <path
           d="m 4273,7867 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5576" />
        <path
           d="m 4334,8295 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5578" />
        <path
           d="m 4394,8723 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5580" />
        <path
           d="m 4454,9151 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5582" />
        <path
           d="m 4492,6246 1,5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5584" />
        <path
           d="m 4909,9210 2,18"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5586" />
        <path
           d="m 4608,7071 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5588" />
        <path
           d="m 4668,7499 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5590" />
        <path
           d="m 4729,7927 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5592" />
        <path
           d="m 4789,8354 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5594" />
        <path
           d="m 4849,8782 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5596" />
        <path
           d="m 4883,5847 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5598" />
        <path
           d="m 5307,8867 2,10"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5600" />
        <path
           d="m 4943,6275 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5602" />
        <path
           d="m 5003,6703 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5604" />
        <path
           d="m 5063,7131 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5606" />
        <path
           d="m 5123,7558 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5608" />
        <path
           d="m 5184,7986 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5610" />
        <path
           d="m 5278,5479 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5612" />
        <path
           d="m 5338,5907 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5614" />
        <path
           d="m 5398,6334 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5616" />
        <path
           d="m 5458,6762 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5618" />
        <path
           d="m 5518,7190 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5620" />
        <path
           d="m 5579,7618 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5622" />
        <path
           d="m 5639,8046 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5624" />
        <path
           d="m 5733,5538 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5626" />
        <path
           d="m 5793,5966 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5628" />
        <path
           d="m 5853,6394 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5630" />
        <path
           d="m 5913,6822 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5632" />
        <path
           d="m 6034,7677 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5634" />
        <path
           d="m 6188,5598 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5636" />
        <path
           d="m 6248,6026 5,35"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5638" />
        <path
           d="m 6368,6881 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5640" />
        <path
           d="m 6643,5657 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5642" />
        <path
           d="m 6703,6085 5,36"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5644" />
        <path
           d="m 7098,5717 5,36 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5646" />
        <path
           d="m 6648,5693 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5648" />
        <path
           d="m 6193,5634 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5650" />
        <path
           d="m 5738,5574 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5652" />
        <path
           d="m 5283,5515 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5654" />
        <path
           d="m 6708,6121 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5656" />
        <path
           d="m 6253,6061 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5658" />
        <path
           d="m 5798,6002 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5660" />
        <path
           d="m 5343,5942 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5662" />
        <path
           d="m 4888,5883 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5664" />
        <path
           d="m 5858,6430 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5666" />
        <path
           d="m 5403,6370 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5668" />
        <path
           d="m 4948,6311 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5670" />
        <path
           d="m 4493,6251 h -3"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5672" />
        <path
           d="m 6373,6917 -37,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5674" />
        <path
           d="m 4519,6674 h -4"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5676" />
        <path
           d="m 5918,6857 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5678" />
        <path
           d="m 5463,6798 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5680" />
        <path
           d="m 5008,6738 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5682" />
        <path
           d="m 4156,7047 -36,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5684" />
        <path
           d="m 5523,7226 -37,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5686" />
        <path
           d="m 5068,7166 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5688" />
        <path
           d="m 4613,7107 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5690" />
        <path
           d="m 6039,7713 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5692" />
        <path
           d="m 5584,7654 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5694" />
        <path
           d="m 5128,7594 -37,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5696" />
        <path
           d="m 4673,7535 -37,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5698" />
        <path
           d="m 4218,7475 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5700" />
        <path
           d="m 5644,8081 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5702" />
        <path
           d="m 5189,8022 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5704" />
        <path
           d="m 4734,7962 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5706" />
        <path
           d="m 4278,7903 -37,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5708" />
        <path
           d="m 5677,8506 -11,-2"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5710" />
        <path
           d="m 4794,8390 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5712" />
        <path
           d="m 4339,8331 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5714" />
        <path
           d="m 3884,8271 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5716" />
        <path
           d="m 5309,8877 h -7"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5718" />
        <path
           d="m 4854,8818 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5720" />
        <path
           d="m 4399,8758 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5722" />
        <path
           d="m 3944,8699 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5724" />
        <path
           d="m 3489,8639 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5726" />
        <path
           d="m 3094,9008 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5728" />
        <path
           d="m 4459,9186 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5730" />
        <path
           d="m 4004,9127 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5732" />
        <path
           d="m 3549,9067 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5734" />
        <path
           d="m 4064,9555 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5736" />
        <path
           d="m 3609,9495 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5738" />
        <path
           d="m 4579,10042 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5740" />
        <path
           d="m 4124,9982 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5742" />
        <path
           d="m 3669,9923 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5744" />
        <path
           d="m 3214,9863 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5746" />
        <path
           d="m 2759,9804 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5748" />
        <path
           d="m 4639,10470 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5750" />
        <path
           d="m 4184,10410 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5752" />
        <path
           d="m 3729,10351 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5754" />
        <path
           d="m 3274,10291 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5756" />
        <path
           d="m 2819,10232 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5758" />
        <path
           d="m 4244,10838 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5760" />
        <path
           d="m 3789,10778 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5762" />
        <path
           d="m 3334,10719 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5764" />
        <path
           d="m 2879,10659 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5766" />
        <path
           d="m 2424,10600 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5768" />
        <path
           d="m 3849,11206 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5770" />
        <path
           d="m 3394,11147 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5772" />
        <path
           d="m 2939,11087 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5774" />
        <path
           d="m 2484,11028 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5776" />
        <path
           d="m 2029,10968 -16,-2"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5778" />
        <path
           d="m 3909,11634 -37,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5780" />
        <path
           d="m 3454,11575 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5782" />
        <path
           d="m 2999,11515 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5784" />
        <path
           d="m 2544,11455 -38,-4"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5786" />
        <path
           d="m 2089,11396 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5788" />
        <path
           d="m 3515,12002 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5790" />
        <path
           d="m 3059,11943 -37,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5792" />
        <path
           d="m 2604,11883 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5794" />
        <path
           d="m 2149,11824 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5796" />
        <path
           d="m 1694,11764 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5798" />
        <path
           d="m 3575,12430 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5800" />
        <path
           d="m 3120,12371 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5802" />
        <path
           d="m 2665,12311 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5804" />
        <path
           d="m 2209,12252 -37,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5806" />
        <path
           d="m 1754,12192 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5808" />
        <path
           d="m 3180,12798 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5810" />
        <path
           d="m 2725,12739 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5812" />
        <path
           d="m 2270,12679 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5814" />
        <path
           d="m 1815,12620 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5816" />
        <path
           d="m 1359,12560 -37,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5818" />
        <path
           d="m 2785,13167 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5820" />
        <path
           d="m 2330,13107 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5822" />
        <path
           d="m 1875,13048 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5824" />
        <path
           d="m 1420,12988 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5826" />
        <path
           d="m 2845,13595 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5828" />
        <path
           d="m 2390,13535 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5830" />
        <path
           d="m 1935,13476 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5832" />
        <path
           d="m 1480,13416 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5834" />
        <path
           d="m 1025,13356 -38,-4"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5836" />
        <path
           d="m 2450,13963 h -1"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5838" />
        <path
           d="m 1995,13903 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5840" />
        <path
           d="m 1540,13844 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5842" />
        <path
           d="m 1085,13784 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5844" />
        <path
           d="m 630,13725 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5846" />
        <path
           d="m 1600,14272 -38,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5848" />
        <path
           d="m 5173,5163 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5850" />
        <path
           d="m 5356,5244 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5852" />
        <path
           d="m 5005,5418 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5854" />
        <path
           d="m 5538,5325 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5856" />
        <path
           d="m 5188,5499 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5858" />
        <path
           d="m 4828,5679 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5860" />
        <path
           d="m 5721,5406 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5862" />
        <path
           d="m 5371,5580 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5864" />
        <path
           d="m 5011,5760 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5866" />
        <path
           d="m 4655,5937 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5868" />
        <path
           d="m 5904,5487 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5870" />
        <path
           d="m 5554,5661 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5872" />
        <path
           d="m 5194,5841 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5874" />
        <path
           d="m 6442,5390 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5876" />
        <path
           d="m 6087,5568 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5878" />
        <path
           d="m 5736,5742 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5880" />
        <path
           d="m 5377,5922 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5882" />
        <path
           d="m 5021,6099 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5884" />
        <path
           d="m 6625,5471 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5886" />
        <path
           d="m 6269,5649 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5888" />
        <path
           d="m 5919,5823 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5890" />
        <path
           d="m 5559,6003 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5892" />
        <path
           d="m 5204,6180 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5894" />
        <path
           d="m 4853,6354 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5896" />
        <path
           d="m 6808,5552 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5898" />
        <path
           d="m 6452,5730 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5900" />
        <path
           d="m 3424,12747 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5902" />
        <path
           d="m 750,13908 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5904" />
        <path
           d="m 1110,13728 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5906" />
        <path
           d="m 1460,13554 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5908" />
        <path
           d="m 1816,13376 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5910" />
        <path
           d="m 2176,13197 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5912" />
        <path
           d="m 2526,13022 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5914" />
        <path
           d="m 2882,12845 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5916" />
        <path
           d="m 3241,12666 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5918" />
        <path
           d="m 568,13827 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5920" />
        <path
           d="m 927,13647 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5922" />
        <path
           d="m 1277,13473 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5924" />
        <path
           d="m 1633,13295 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5926" />
        <path
           d="m 1993,13116 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5928" />
        <path
           d="m 2343,12941 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5930" />
        <path
           d="m 2699,12764 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5932" />
        <path
           d="m 3059,12585 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5934" />
        <path
           d="m 3409,12410 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5936" />
        <path
           d="m 745,13566 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5938" />
        <path
           d="m 1095,13392 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5940" />
        <path
           d="m 1450,13214 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5942" />
        <path
           d="m 1810,13035 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5944" />
        <path
           d="m 2160,12860 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5946" />
        <path
           d="m 2516,12683 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5948" />
        <path
           d="m 2876,12504 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5950" />
        <path
           d="m 3226,12329 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5952" />
        <path
           d="m 3582,12152 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5954" />
        <path
           d="m 912,13311 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5956" />
        <path
           d="m 1268,13133 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5958" />
        <path
           d="m 1627,12954 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5960" />
        <path
           d="m 1978,12779 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5962" />
        <path
           d="m 2333,12602 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5964" />
        <path
           d="m 2693,12423 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5966" />
        <path
           d="m 3043,12248 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5968" />
        <path
           d="m 3399,12071 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5970" />
        <path
           d="m 3759,11891 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5972" />
        <path
           d="m 1085,13052 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5974" />
        <path
           d="m 1445,12873 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5976" />
        <path
           d="m 1795,12698 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5978" />
        <path
           d="m 2151,12521 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5980" />
        <path
           d="m 2510,12342 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5982" />
        <path
           d="m 2861,12167 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5984" />
        <path
           d="m 3216,11990 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5986" />
        <path
           d="m 3576,11810 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5988" />
        <path
           d="m 3926,11636 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5990" />
        <path
           d="m 1262,12792 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5992" />
        <path
           d="m 1612,12617 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5994" />
        <path
           d="m 1968,12440 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5996" />
        <path
           d="m 2328,12261 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path5998" />
        <path
           d="m 2678,12086 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6000" />
        <path
           d="m 3034,11909 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6002" />
        <path
           d="m 3393,11729 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6004" />
        <path
           d="m 3743,11555 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6006" />
        <path
           d="m 4099,11377 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6008" />
        <path
           d="m 1429,12536 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6010" />
        <path
           d="m 1785,12359 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6012" />
        <path
           d="m 2145,12180 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6014" />
        <path
           d="m 2495,12005 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6016" />
        <path
           d="m 2851,11828 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6018" />
        <path
           d="m 3211,11648 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6020" />
        <path
           d="m 3561,11474 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6022" />
        <path
           d="m 3916,11296 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6024" />
        <path
           d="m 4276,11117 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6026" />
        <path
           d="m 1247,12455 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6028" />
        <path
           d="m 1602,12278 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6030" />
        <path
           d="m 1962,12099 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6032" />
        <path
           d="m 2312,11924 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6034" />
        <path
           d="m 2668,11747 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6036" />
        <path
           d="m 3028,11567 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6038" />
        <path
           d="m 3378,11393 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6040" />
        <path
           d="m 3734,11215 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6042" />
        <path
           d="m 4093,11036 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6044" />
        <path
           d="m 1420,12197 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6046" />
        <path
           d="m 1779,12018 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6048" />
        <path
           d="m 2130,11843 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6050" />
        <path
           d="m 2485,11666 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6052" />
        <path
           d="m 2845,11486 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6054" />
        <path
           d="m 3195,11312 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6056" />
        <path
           d="m 3551,11134 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6058" />
        <path
           d="m 3911,10955 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6060" />
        <path
           d="m 1597,11937 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6062" />
        <path
           d="m 1947,11762 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6064" />
        <path
           d="m 2303,11585 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6066" />
        <path
           d="m 2662,11405 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6068" />
        <path
           d="m 3013,11231 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6070" />
        <path
           d="m 3368,11053 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6072" />
        <path
           d="m 3728,10874 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6074" />
        <path
           d="m 4434,10522 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6076" />
        <path
           d="m 1764,11681 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6078" />
        <path
           d="m 2120,11504 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6080" />
        <path
           d="m 2480,11324 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6082" />
        <path
           d="m 2830,11150 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6084" />
        <path
           d="m 3186,10972 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6086" />
        <path
           d="m 3545,10793 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6088" />
        <path
           d="m 3895,10619 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6090" />
        <path
           d="m 4251,10441 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6092" />
        <path
           d="m 4611,10262 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6094" />
        <path
           d="m 1937,11423 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6096" />
        <path
           d="m 2297,11243 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6098" />
        <path
           d="m 2647,11069 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6100" />
        <path
           d="m 3003,10891 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6102" />
        <path
           d="m 3363,10712 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6104" />
        <path
           d="m 3713,10538 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6106" />
        <path
           d="m 4068,10360 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6108" />
        <path
           d="m 4428,10181 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6110" />
        <path
           d="m 4778,10006 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6112" />
        <path
           d="m 2114,11162 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6114" />
        <path
           d="m 2464,10988 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6116" />
        <path
           d="m 2820,10810 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6118" />
        <path
           d="m 3180,10631 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6120" />
        <path
           d="m 3530,10457 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6122" />
        <path
           d="m 3886,10279 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6124" />
        <path
           d="m 4245,10100 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6126" />
        <path
           d="m 4596,9925 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6128" />
        <path
           d="m 2282,10907 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6130" />
        <path
           d="m 2637,10729 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6132" />
        <path
           d="m 2997,10550 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6134" />
        <path
           d="m 3347,10376 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6136" />
        <path
           d="m 3703,10198 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6138" />
        <path
           d="m 4063,10019 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6140" />
        <path
           d="m 4413,9844 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6142" />
        <path
           d="m 2099,10826 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6144" />
        <path
           d="m 2455,10648 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6146" />
        <path
           d="m 2814,10469 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6148" />
        <path
           d="m 3165,10295 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6150" />
        <path
           d="m 3520,10117 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6152" />
        <path
           d="m 3880,9938 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6154" />
        <path
           d="m 4230,9763 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6156" />
        <path
           d="m 5296,9232 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6158" />
        <path
           d="m 2272,10567 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6160" />
        <path
           d="m 2632,10388 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6162" />
        <path
           d="m 2982,10214 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6164" />
        <path
           d="m 3338,10036 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6166" />
        <path
           d="m 3697,9857 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6168" />
        <path
           d="m 4047,9682 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6170" />
        <path
           d="m 4403,9505 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6172" />
        <path
           d="m 2449,10307 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6174" />
        <path
           d="m 2799,10133 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6176" />
        <path
           d="m 3155,9955 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6178" />
        <path
           d="m 3515,9776 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6180" />
        <path
           d="m 3865,9601 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6182" />
        <path
           d="m 4220,9424 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6184" />
        <path
           d="m 4580,9244 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6186" />
        <path
           d="m 3332,9695 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6188" />
        <path
           d="m 3682,9520 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6190" />
        <path
           d="m 4038,9343 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6192" />
        <path
           d="m 4397,9163 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6194" />
        <path
           d="m 4748,8989 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6196" />
        <path
           d="m 2616,10052 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6198" />
        <path
           d="m 5463,8632 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6200" />
        <path
           d="m 3149,9614 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6202" />
        <path
           d="m 3499,9439 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6204" />
        <path
           d="m 3855,9262 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6206" />
        <path
           d="m 4215,9082 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6208" />
        <path
           d="m 4565,8908 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6210" />
        <path
           d="m 4921,8731 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6212" />
        <path
           d="m 5630,8377 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6214" />
        <path
           d="m 3317,9358 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6216" />
        <path
           d="m 3672,9181 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6218" />
        <path
           d="m 4032,9001 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6220" />
        <path
           d="m 4382,8827 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6222" />
        <path
           d="m 4738,8650 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6224" />
        <path
           d="m 5098,8470 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6226" />
        <path
           d="m 2966,9533 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6228" />
        <path
           d="m 5448,8296 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6230" />
        <path
           d="m 5804,8118 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6232" />
        <path
           d="m 3490,9100 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6234" />
        <path
           d="m 3849,8920 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6236" />
        <path
           d="m 4199,8746 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6238" />
        <path
           d="m 4555,8569 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6240" />
        <path
           d="m 4915,8389 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6242" />
        <path
           d="m 5265,8215 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6244" />
        <path
           d="m 5621,8037 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6246" />
        <path
           d="m 5981,7858 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6248" />
        <path
           d="m 2951,9196 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6250" />
        <path
           d="m 3667,8839 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6252" />
        <path
           d="m 4017,8665 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6254" />
        <path
           d="m 4372,8488 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6256" />
        <path
           d="m 4732,8308 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6258" />
        <path
           d="m 5082,8134 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6260" />
        <path
           d="m 5438,7956 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6262" />
        <path
           d="m 5798,7777 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6264" />
        <path
           d="m 6148,7602 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6266" />
        <path
           d="m 3484,8758 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6268" />
        <path
           d="m 3834,8584 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6270" />
        <path
           d="m 4190,8407 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6272" />
        <path
           d="m 4549,8227 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6274" />
        <path
           d="m 4900,8053 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6276" />
        <path
           d="m 5255,7875 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6278" />
        <path
           d="m 5615,7696 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6280" />
        <path
           d="m 3124,8938 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6282" />
        <path
           d="m 3301,8677 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6284" />
        <path
           d="m 3651,8503 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6286" />
        <path
           d="m 4007,8326 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6288" />
        <path
           d="m 4367,8146 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6290" />
        <path
           d="m 4717,7972 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6292" />
        <path
           d="m 5073,7794 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6294" />
        <path
           d="m 5432,7615 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6296" />
        <path
           d="m 3824,8245 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6298" />
        <path
           d="m 4184,8065 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6300" />
        <path
           d="m 4534,7891 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6302" />
        <path
           d="m 4890,7713 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6304" />
        <path
           d="m 5250,7534 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6306" />
        <path
           d="m 5600,7359 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6308" />
        <path
           d="m 6315,7003 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6310" />
        <path
           d="m 4001,7984 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6312" />
        <path
           d="m 4351,7810 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6314" />
        <path
           d="m 4707,7632 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6316" />
        <path
           d="m 5067,7453 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6318" />
        <path
           d="m 5417,7278 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6320" />
        <path
           d="m 5773,7101 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6322" />
        <path
           d="m 4169,7729 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6324" />
        <path
           d="m 4524,7551 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6326" />
        <path
           d="m 4884,7372 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6328" />
        <path
           d="m 5234,7197 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6330" />
        <path
           d="m 5590,7020 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6332" />
        <path
           d="m 5950,6841 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6334" />
        <path
           d="m 3986,7648 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6336" />
        <path
           d="m 4342,7470 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6338" />
        <path
           d="m 4701,7291 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6340" />
        <path
           d="m 5052,7116 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6342" />
        <path
           d="m 5407,6939 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6344" />
        <path
           d="m 5767,6760 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6346" />
        <path
           d="m 6833,6228 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6348" />
        <path
           d="m 3803,7567 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6350" />
        <path
           d="m 4159,7389 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6352" />
        <path
           d="m 4519,7210 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6354" />
        <path
           d="m 4869,7035 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6356" />
        <path
           d="m 5225,6858 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6358" />
        <path
           d="m 5584,6679 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6360" />
        <path
           d="m 5935,6504 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6362" />
        <path
           d="m 6650,6147 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6364" />
        <path
           d="m 7000,5973 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6366" />
        <path
           d="m 4686,6954 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6368" />
        <path
           d="m 5042,6777 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6370" />
        <path
           d="m 5402,6598 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6372" />
        <path
           d="m 5752,6423 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6374" />
        <path
           d="m 6108,6246 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6376" />
        <path
           d="m 3976,7308 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6378" />
        <path
           d="m 6467,6066 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6380" />
        <path
           d="m 6817,5892 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6382" />
        <path
           d="m 4153,7048 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6384" />
        <path
           d="m 4503,6873 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6386" />
        <path
           d="m 4859,6696 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6388" />
        <path
           d="m 5219,6516 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6390" />
        <path
           d="m 5569,6342 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6392" />
        <path
           d="m 5925,6165 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6394" />
        <path
           d="m 6285,5985 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6396" />
        <path
           d="m 6635,5811 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6398" />
        <path
           d="m 6990,5633 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6400" />
        <path
           d="m 4321,6792 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6402" />
        <path
           d="m 4676,6615 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6404" />
        <path
           d="m 5036,6435 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6406" />
        <path
           d="m 5386,6261 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6408" />
        <path
           d="m 5742,6084 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6410" />
        <path
           d="m 6102,5904 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6412" />
        <path
           d="m 6917,5749 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6414" />
        <path
           d="m 1161,14058 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6416" />
        <path
           d="m 1372,13739 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6418" />
        <path
           d="m 1499,13548 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6420" />
        <path
           d="m 1582,13421 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6422" />
        <path
           d="m 1793,13103 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6424" />
        <path
           d="m 1920,12912 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6426" />
        <path
           d="m 2003,12785 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6428" />
        <path
           d="m 2214,12467 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6430" />
        <path
           d="m 2341,12275 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6432" />
        <path
           d="m 2424,12149 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6434" />
        <path
           d="m 2635,11830 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6436" />
        <path
           d="m 2762,11639 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6438" />
        <path
           d="m 2845,11513 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6440" />
        <path
           d="m 3056,11194 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6442" />
        <path
           d="m 3183,11003 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6444" />
        <path
           d="m 3266,10877 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6446" />
        <path
           d="m 3477,10558 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6448" />
        <path
           d="m 3604,10367 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6450" />
        <path
           d="m 3688,10241 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6452" />
        <path
           d="m 3899,9922 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6454" />
        <path
           d="m 4025,9731 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6456" />
        <path
           d="m 4109,9604 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6458" />
        <path
           d="m 4320,9286 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6460" />
        <path
           d="m 4446,9094 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6462" />
        <path
           d="m 4530,8968 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6464" />
        <path
           d="m 4741,8649 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6466" />
        <path
           d="m 4867,8458 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6468" />
        <path
           d="m 4951,8332 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6470" />
        <path
           d="m 5162,8013 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6472" />
        <path
           d="m 5288,7822 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6474" />
        <path
           d="m 5372,7696 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6476" />
        <path
           d="m 5583,7377 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6478" />
        <path
           d="m 5709,7186 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6480" />
        <path
           d="m 5793,7060 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6482" />
        <path
           d="m 6004,6741 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6484" />
        <path
           d="m 6425,6105 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6486" />
        <path
           d="m 6552,5914 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6488" />
        <path
           d="m 6635,5787 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6490" />
        <path
           d="m 6846,5468 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6492" />
        <path
           d="m 1090,13777 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6494" />
        <path
           d="m 1217,13586 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6496" />
        <path
           d="m 1300,13460 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6498" />
        <path
           d="m 1511,13141 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6500" />
        <path
           d="m 1638,12950 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6502" />
        <path
           d="m 1721,12823 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6504" />
        <path
           d="m 1932,12505 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6506" />
        <path
           d="m 2059,12314 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6508" />
        <path
           d="m 2142,12187 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6510" />
        <path
           d="m 2353,11869 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6512" />
        <path
           d="m 2480,11677 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6514" />
        <path
           d="m 2563,11551 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6516" />
        <path
           d="m 2774,11232 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6518" />
        <path
           d="m 2901,11041 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6520" />
        <path
           d="m 2985,10915 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6522" />
        <path
           d="m 3196,10596 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6524" />
        <path
           d="m 3322,10405 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6526" />
        <path
           d="m 3406,10279 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6528" />
        <path
           d="m 3617,9960 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6530" />
        <path
           d="m 3743,9769 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6532" />
        <path
           d="m 3827,9642 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6534" />
        <path
           d="m 4038,9324 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6536" />
        <path
           d="m 4164,9133 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6538" />
        <path
           d="m 4248,9006 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6540" />
        <path
           d="m 4459,8688 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6542" />
        <path
           d="m 4585,8496 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6544" />
        <path
           d="m 4669,8370 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6546" />
        <path
           d="m 4880,8051 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6548" />
        <path
           d="m 5006,7860 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6550" />
        <path
           d="m 5090,7734 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6552" />
        <path
           d="m 5301,7415 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6554" />
        <path
           d="m 5427,7224 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6556" />
        <path
           d="m 5511,7098 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6558" />
        <path
           d="m 5722,6779 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6560" />
        <path
           d="m 5849,6588 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6562" />
        <path
           d="m 5932,6462 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6564" />
        <path
           d="m 6143,6143 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6566" />
        <path
           d="m 6270,5952 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6568" />
        <path
           d="m 6353,5825 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6570" />
        <path
           d="m 6564,5507 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6572" />
        <path
           d="m 808,13815 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6574" />
        <path
           d="m 935,13624 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6576" />
        <path
           d="m 1018,13498 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6578" />
        <path
           d="m 1229,13179 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6580" />
        <path
           d="m 1356,12988 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6582" />
        <path
           d="m 1439,12862 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6584" />
        <path
           d="m 1650,12543 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6586" />
        <path
           d="m 1777,12352 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6588" />
        <path
           d="m 1860,12225 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6590" />
        <path
           d="m 2071,11907 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6592" />
        <path
           d="m 2198,11715 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6594" />
        <path
           d="m 2282,11589 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6596" />
        <path
           d="m 2493,11270 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6598" />
        <path
           d="m 2703,10953 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6600" />
        <path
           d="m 2914,10634 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6602" />
        <path
           d="m 3040,10443 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6604" />
        <path
           d="m 3124,10317 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6606" />
        <path
           d="m 3335,9998 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6608" />
        <path
           d="m 3461,9807 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6610" />
        <path
           d="m 3545,9681 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6612" />
        <path
           d="m 3756,9362 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6614" />
        <path
           d="m 3882,9171 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6616" />
        <path
           d="m 3966,9044 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6618" />
        <path
           d="m 4177,8726 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6620" />
        <path
           d="m 4303,8535 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6622" />
        <path
           d="m 4387,8408 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6624" />
        <path
           d="m 4598,8089 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6626" />
        <path
           d="m 4724,7898 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6628" />
        <path
           d="m 4808,7772 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6630" />
        <path
           d="m 5019,7453 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6632" />
        <path
           d="m 5146,7262 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6634" />
        <path
           d="m 5229,7136 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6636" />
        <path
           d="m 5440,6817 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6638" />
        <path
           d="m 5567,6626 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6640" />
        <path
           d="m 5650,6500 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6642" />
        <path
           d="m 5861,6181 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6644" />
        <path
           d="m 5988,5990 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6646" />
        <path
           d="m 6071,5863 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6648" />
        <path
           d="m 6282,5545 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6650" />
        <path
           d="m 653,13662 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6652" />
        <path
           d="m 736,13536 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6654" />
        <path
           d="m 947,13217 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6656" />
        <path
           d="m 1074,13026 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6658" />
        <path
           d="m 1158,12900 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6660" />
        <path
           d="m 1368,12581 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6662" />
        <path
           d="m 1495,12390 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6664" />
        <path
           d="m 1579,12263 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6666" />
        <path
           d="m 1790,11945 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6668" />
        <path
           d="m 1916,11754 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6670" />
        <path
           d="m 2000,11627 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6672" />
        <path
           d="m 2211,11309 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6674" />
        <path
           d="m 2337,11117 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6676" />
        <path
           d="m 2421,10991 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6678" />
        <path
           d="m 2632,10672 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6680" />
        <path
           d="m 2758,10481 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6682" />
        <path
           d="m 2842,10355 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6684" />
        <path
           d="m 3053,10036 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6686" />
        <path
           d="m 3179,9845 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6688" />
        <path
           d="m 3263,9719 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6690" />
        <path
           d="m 3474,9400 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6692" />
        <path
           d="m 3600,9209 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6694" />
        <path
           d="m 3684,9083 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6696" />
        <path
           d="m 3895,8764 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6698" />
        <path
           d="m 4021,8573 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6700" />
        <path
           d="m 4105,8446 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6702" />
        <path
           d="m 4316,8128 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6704" />
        <path
           d="m 4443,7936 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6706" />
        <path
           d="m 4526,7810 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6708" />
        <path
           d="m 4737,7491 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6710" />
        <path
           d="m 4864,7300 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6712" />
        <path
           d="m 4947,7174 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6714" />
        <path
           d="m 5158,6855 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6716" />
        <path
           d="m 5285,6664 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6718" />
        <path
           d="m 5368,6538 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6720" />
        <path
           d="m 5579,6219 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6722" />
        <path
           d="m 5706,6028 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6724" />
        <path
           d="m 5789,5902 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6726" />
        <path
           d="m 6000,5583 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6728" />
        <path
           d="m 6127,5392 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6730" />
        <path
           d="m 3319,9247 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6732" />
        <path
           d="m 1508,11983 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6734" />
        <path
           d="m 1634,11792 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6736" />
        <path
           d="m 1718,11665 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6738" />
        <path
           d="m 1929,11347 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6740" />
        <path
           d="m 2055,11156 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6742" />
        <path
           d="m 2139,11029 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6744" />
        <path
           d="m 2350,10711 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6746" />
        <path
           d="m 2476,10519 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6748" />
        <path
           d="m 2560,10393 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6750" />
        <path
           d="m 2771,10074 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6752" />
        <path
           d="m 2897,9883 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6754" />
        <path
           d="m 3402,9121 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6756" />
        <path
           d="m 3613,8802 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6758" />
        <path
           d="m 3740,8611 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6760" />
        <path
           d="m 3823,8484 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6762" />
        <path
           d="m 4034,8166 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6764" />
        <path
           d="m 4161,7975 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6766" />
        <path
           d="m 4244,7848 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6768" />
        <path
           d="m 4455,7530 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6770" />
        <path
           d="m 4582,7338 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6772" />
        <path
           d="m 4665,7212 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6774" />
        <path
           d="m 4876,6893 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6776" />
        <path
           d="m 5003,6702 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6778" />
        <path
           d="m 5086,6576 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6780" />
        <path
           d="m 5297,6257 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6782" />
        <path
           d="m 5424,6066 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6784" />
        <path
           d="m 5508,5940 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6786" />
        <path
           d="m 5719,5621 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6788" />
        <path
           d="m 5845,5430 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6790" />
        <path
           d="m 5929,5304 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6792" />
        <path
           d="m 3458,8649 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6794" />
        <path
           d="m 3541,8523 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6796" />
        <path
           d="m 3331,8840 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6798" />
        <path
           d="m 4173,7568 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6800" />
        <path
           d="m 3120,9159 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6802" />
        <path
           d="m 4300,7377 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6804" />
        <path
           d="m 2489,10112 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6806" />
        <path
           d="m 2616,9921 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6808" />
        <path
           d="m 2699,9795 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6810" />
        <path
           d="m 2910,9476 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6812" />
        <path
           d="m 4594,6931 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6814" />
        <path
           d="m 4721,6740 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6816" />
        <path
           d="m 4805,6614 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6818" />
        <path
           d="m 5016,6295 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6820" />
        <path
           d="m 5142,6104 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6822" />
        <path
           d="m 5226,5978 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6824" />
        <path
           d="m 5437,5659 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6826" />
        <path
           d="m 5563,5468 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6828" />
        <path
           d="m 5647,5342 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6830" />
        <path
           d="m 3891,7606 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6832" />
        <path
           d="m 4018,7415 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6834" />
        <path
           d="m 4102,7288 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6836" />
        <path
           d="m 3470,8242 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6838" />
        <path
           d="m 3597,8051 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6840" />
        <path
           d="m 3680,7925 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6842" />
        <path
           d="m 4439,6778 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6844" />
        <path
           d="m 5155,5697 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6846" />
        <path
           d="m 5281,5506 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6848" />
        <path
           d="m 5365,5380 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6850" />
        <path
           d="m 4873,5735 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6852" />
        <path
           d="m 4999,5544 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6854" />
        <path
           d="m 5083,5418 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6856" />
        <path
           d="m 4452,6372 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6858" />
        <path
           d="m 4578,6180 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6860" />
        <path
           d="m 4662,6054 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6862" />
        <path
           d="m 2395,14637 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6864" />
        <path
           d="m 2212,14556 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6866" />
        <path
           d="m 2029,14475 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6868" />
        <path
           d="m 1847,14394 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6870" />
        <path
           d="m 1664,14313 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6872" />
        <path
           d="m 2024,14133 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6874" />
        <path
           d="m 2730,13781 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6876" />
        <path
           d="m 1481,14232 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6878" />
        <path
           d="m 1841,14052 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6880" />
        <path
           d="m 2547,13700 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6882" />
        <path
           d="m 2907,13521 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6884" />
        <path
           d="m 1298,14151 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6886" />
        <path
           d="m 1658,13971 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6888" />
        <path
           d="m 2008,13797 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6890" />
        <path
           d="m 2364,13619 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6892" />
        <path
           d="m 2724,13440 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6894" />
        <path
           d="m 3074,13265 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6896" />
        <path
           d="m 1116,14070 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6898" />
        <path
           d="m 1475,13890 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6900" />
        <path
           d="m 1826,13716 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6902" />
        <path
           d="m 2181,13538 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6904" />
        <path
           d="m 2541,13359 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6906" />
        <path
           d="m 2891,13184 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6908" />
        <path
           d="m 3247,13007 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6910" />
        <path
           d="m 933,13989 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6912" />
        <path
           d="m 1293,13809 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6914" />
        <path
           d="m 1643,13635 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6916" />
        <path
           d="m 1999,13457 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6918" />
        <path
           d="m 2358,13278 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6920" />
        <path
           d="m 2709,13103 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6922" />
        <path
           d="m 3064,12926 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6924" />
        <path
           d="m 3633,11380 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6926" />
        <path
           d="m 3580,10915 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6928" />
        <path
           d="m 3563,10766 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6930" />
        <path
           d="m 3493,10149 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6932" />
        <path
           d="m 3440,9684 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6934" />
        <path
           d="m 3423,9535 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6936" />
        <path
           d="m 3224,9212 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6938" />
        <path
           d="m 3592,12440 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6940" />
        <path
           d="m 3575,12291 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6942" />
        <path
           d="m 3505,11674 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6944" />
        <path
           d="m 3452,11209 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6946" />
        <path
           d="m 3435,11060 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6948" />
        <path
           d="m 3365,10443 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6950" />
        <path
           d="m 3312,9978 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6952" />
        <path
           d="m 3295,9829 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6954" />
        <path
           d="m 3447,12585 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6956" />
        <path
           d="m 3377,11968 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6958" />
        <path
           d="m 3324,11503 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6960" />
        <path
           d="m 3307,11354 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6962" />
        <path
           d="m 3236,10737 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6964" />
        <path
           d="m 3183,10272 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6966" />
        <path
           d="m 3166,10123 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6968" />
        <path
           d="m 3043,9041 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6970" />
        <path
           d="m 3319,12879 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6972" />
        <path
           d="m 3248,12261 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6974" />
        <path
           d="m 3195,11796 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6976" />
        <path
           d="m 3178,11647 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6978" />
        <path
           d="m 3108,11030 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6980" />
        <path
           d="m 3055,10565 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6982" />
        <path
           d="m 3038,10416 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6984" />
        <path
           d="m 2915,9334 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6986" />
        <path
           d="m 3190,13172 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6988" />
        <path
           d="m 3120,12555 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6990" />
        <path
           d="m 3067,12090 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6992" />
        <path
           d="m 3050,11941 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6994" />
        <path
           d="m 2980,11324 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6996" />
        <path
           d="m 2927,10859 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path6998" />
        <path
           d="m 2910,10710 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7000" />
        <path
           d="m 2840,10093 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7002" />
        <path
           d="m 2787,9628 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7004" />
        <path
           d="m 3062,13466 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7006" />
        <path
           d="m 2992,12849 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7008" />
        <path
           d="m 2939,12384 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7010" />
        <path
           d="m 2922,12235 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7012" />
        <path
           d="m 2852,11618 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7014" />
        <path
           d="m 2799,11153 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7016" />
        <path
           d="m 2782,11004 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7018" />
        <path
           d="m 2711,10387 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7020" />
        <path
           d="m 2658,9922 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7022" />
        <path
           d="m 2641,9773 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7024" />
        <path
           d="m 2864,13143 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7026" />
        <path
           d="m 2811,12678 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7028" />
        <path
           d="m 2794,12529 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7030" />
        <path
           d="m 2723,11912 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7032" />
        <path
           d="m 2670,11447 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7034" />
        <path
           d="m 2653,11298 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7036" />
        <path
           d="m 2583,10681 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7038" />
        <path
           d="m 2530,10216 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7040" />
        <path
           d="m 2513,10067 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7042" />
        <path
           d="m 2735,13437 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7044" />
        <path
           d="m 2682,12972 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7046" />
        <path
           d="m 2665,12823 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7048" />
        <path
           d="m 2595,12206 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7050" />
        <path
           d="m 2542,11741 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7052" />
        <path
           d="m 2525,11592 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7054" />
        <path
           d="m 2455,10975 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7056" />
        <path
           d="m 2402,10510 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7058" />
        <path
           d="m 2385,10361 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7060" />
        <path
           d="m 2607,13731 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7062" />
        <path
           d="m 2554,13266 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7064" />
        <path
           d="m 2537,13117 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7066" />
        <path
           d="m 2467,12500 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7068" />
        <path
           d="m 2414,12035 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7070" />
        <path
           d="m 2397,11885 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7072" />
        <path
           d="m 2327,11268 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7074" />
        <path
           d="m 2274,10803 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7076" />
        <path
           d="m 2257,10654 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7078" />
        <path
           d="m 2426,13559 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7080" />
        <path
           d="m 2409,13410 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7082" />
        <path
           d="m 2339,12793 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7084" />
        <path
           d="m 2286,12328 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7086" />
        <path
           d="m 2269,12179 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7088" />
        <path
           d="m 2198,11562 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7090" />
        <path
           d="m 2145,11097 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7092" />
        <path
           d="m 2128,10948 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7094" />
        <path
           d="m 2298,13853 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7096" />
        <path
           d="m 2281,13704 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7098" />
        <path
           d="m 2210,13087 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7100" />
        <path
           d="m 2157,12622 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7102" />
        <path
           d="m 2140,12473 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7104" />
        <path
           d="m 2070,11856 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7106" />
        <path
           d="m 2017,11391 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7108" />
        <path
           d="m 2000,11242 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7110" />
        <path
           d="m 2222,14612 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7112" />
        <path
           d="m 2082,13381 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7114" />
        <path
           d="m 2029,12916 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7116" />
        <path
           d="m 2012,12767 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7118" />
        <path
           d="m 1942,12150 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7120" />
        <path
           d="m 1889,11685 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7122" />
        <path
           d="m 1872,11536 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7124" />
        <path
           d="m 2041,14441 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7126" />
        <path
           d="m 1954,13675 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7128" />
        <path
           d="m 1901,13210 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7130" />
        <path
           d="m 1884,13061 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7132" />
        <path
           d="m 1814,12444 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7134" />
        <path
           d="m 1761,11979 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7136" />
        <path
           d="m 1744,11830 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7138" />
        <path
           d="m 1826,13969 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7140" />
        <path
           d="m 1773,13504 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7142" />
        <path
           d="m 1756,13355 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7144" />
        <path
           d="m 1685,12738 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7146" />
        <path
           d="m 1632,12273 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7148" />
        <path
           d="m 1615,12123 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7150" />
        <path
           d="m 1697,14262 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7152" />
        <path
           d="m 1644,13797 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7154" />
        <path
           d="m 1627,13648 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7156" />
        <path
           d="m 1557,13031 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7158" />
        <path
           d="m 1504,12566 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7160" />
        <path
           d="m 1487,12417 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7162" />
        <path
           d="m 1516,14091 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7164" />
        <path
           d="m 1499,13942 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7166" />
        <path
           d="m 1429,13325 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7168" />
        <path
           d="m 1376,12860 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7170" />
        <path
           d="m 1359,12711 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7172" />
        <path
           d="m 1371,14236 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7174" />
        <path
           d="m 1301,13619 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7176" />
        <path
           d="m 1248,13154 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7178" />
        <path
           d="m 1231,13005 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7180" />
        <path
           d="m 1172,13913 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7182" />
        <path
           d="m 1119,13448 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7184" />
        <path
           d="m 1102,13299 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7186" />
        <path
           d="m 991,13742 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7188" />
        <path
           d="m 974,13593 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7190" />
        <path
           d="m 846,13886 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7192" />
        <path
           d="m 2348,14591 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7194" />
        <path
           d="m 2769,13955 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7196" />
        <path
           d="m 2852,13829 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7198" />
        <path
           d="m 2149,14503 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7200" />
        <path
           d="m 2571,13867 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7202" />
        <path
           d="m 2781,13548 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7204" />
        <path
           d="m 2908,13357 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7206" />
        <path
           d="m 2992,13231 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7208" />
        <path
           d="m 3203,12912 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7210" />
        <path
           d="m 3329,12721 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7212" />
        <path
           d="m 3413,12595 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7214" />
        <path
           d="m 3624,12276 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7216" />
        <path
           d="m 3750,12085 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7218" />
        <path
           d="m 3834,11958 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7220" />
        <path
           d="m 2500,13586 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7222" />
        <path
           d="m 2626,13395 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7224" />
        <path
           d="m 2710,13269 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7226" />
        <path
           d="m 2921,12950 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7228" />
        <path
           d="m 3047,12759 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7230" />
        <path
           d="m 3131,12633 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7232" />
        <path
           d="m 3342,12314 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7234" />
        <path
           d="m 3468,12123 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7236" />
        <path
           d="m 3552,11997 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7238" />
        <path
           d="m 3763,11678 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7240" />
        <path
           d="m 3889,11487 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7242" />
        <path
           d="m 3973,11360 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7244" />
        <path
           d="m 4184,11042 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7246" />
        <path
           d="m 4310,10851 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7248" />
        <path
           d="m 4605,10405 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7250" />
        <path
           d="m 4732,10214 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7252" />
        <path
           d="m 4815,10088 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7254" />
        <path
           d="m 4323,10444 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7256" />
        <path
           d="m 4450,10252 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7258" />
        <path
           d="m 4533,10126 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7260" />
        <path
           d="m 1797,14261 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7262" />
        <path
           d="m 1923,14070 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7264" />
        <path
           d="m 2007,13943 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7266" />
        <path
           d="m 2218,13625 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7268" />
        <path
           d="m 2344,13433 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7270" />
        <path
           d="m 2428,13307 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7272" />
        <path
           d="m 2639,12988 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7274" />
        <path
           d="m 2765,12797 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7276" />
        <path
           d="m 2849,12671 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7278" />
        <path
           d="m 3060,12352 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7280" />
        <path
           d="m 3186,12161 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7282" />
        <path
           d="m 3270,12035 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7284" />
        <path
           d="m 3481,11716 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7286" />
        <path
           d="m 3607,11525 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7288" />
        <path
           d="m 3691,11399 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7290" />
        <path
           d="m 3902,11080 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7292" />
        <path
           d="m 4029,10889 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7294" />
        <path
           d="m 4112,10762 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7296" />
        <path
           d="m 5165,9171 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7298" />
        <path
           d="m 5292,8980 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7300" />
        <path
           d="m 5375,8854 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7302" />
        <path
           d="m 5586,8535 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7304" />
        <path
           d="m 5713,8344 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7306" />
        <path
           d="m 5797,8218 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7308" />
        <path
           d="m 5431,8382 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7310" />
        <path
           d="m 5515,8256 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7312" />
        <path
           d="m 5726,7937 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7314" />
        <path
           d="m 5852,7746 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7316" />
        <path
           d="m 4883,9209 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7318" />
        <path
           d="m 6147,7301 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7320" />
        <path
           d="m 6273,7110 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7322" />
        <path
           d="m 6357,6983 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7324" />
        <path
           d="m 1515,14299 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7326" />
        <path
           d="m 1641,14108 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7328" />
        <path
           d="m 1725,13981 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7330" />
        <path
           d="m 1936,13663 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7332" />
        <path
           d="m 2062,13472 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7334" />
        <path
           d="m 2146,13345 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7336" />
        <path
           d="m 2357,13026 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7338" />
        <path
           d="m 2483,12835 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7340" />
        <path
           d="m 2567,12709 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7342" />
        <path
           d="m 2778,12390 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7344" />
        <path
           d="m 2904,12199 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7346" />
        <path
           d="m 2988,12073 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7348" />
        <path
           d="m 3199,11754 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7350" />
        <path
           d="m 3326,11563 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7352" />
        <path
           d="m 3409,11437 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7354" />
        <path
           d="m 3620,11118 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7356" />
        <path
           d="m 3747,10927 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7358" />
        <path
           d="m 3830,10800 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7360" />
        <path
           d="m 4041,10482 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7362" />
        <path
           d="m 4168,10291 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7364" />
        <path
           d="m 4251,10164 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7366" />
        <path
           d="m 4462,9846 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7368" />
        <path
           d="m 4728,9056 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7370" />
        <path
           d="m 4812,8930 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7372" />
        <path
           d="m 5023,8611 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7374" />
        <path
           d="m 5149,8420 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7376" />
        <path
           d="m 5233,8294 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7378" />
        <path
           d="m 5444,7975 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7380" />
        <path
           d="m 5570,7784 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7382" />
        <path
           d="m 5654,7658 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7384" />
        <path
           d="m 1359,14146 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7386" />
        <path
           d="m 1443,14020 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7388" />
        <path
           d="m 1654,13701 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7390" />
        <path
           d="m 1780,13510 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7392" />
        <path
           d="m 1864,13383 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7394" />
        <path
           d="m 2075,13065 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7396" />
        <path
           d="m 2201,12873 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7398" />
        <path
           d="m 2285,12747 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7400" />
        <path
           d="m 2496,12428 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7402" />
        <path
           d="m 2623,12237 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7404" />
        <path
           d="m 2706,12111 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7406" />
        <path
           d="m 2917,11792 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7408" />
        <path
           d="m 3044,11601 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7410" />
        <path
           d="m 3127,11475 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7412" />
        <path
           d="m 3338,11156 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7414" />
        <path
           d="m 3465,10965 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7416" />
        <path
           d="m 3548,10839 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7418" />
        <path
           d="m 3759,10520 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7420" />
        <path
           d="m 3886,10329 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7422" />
        <path
           d="m 3969,10202 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7424" />
        <path
           d="m 4180,9884 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7426" />
        <path
           d="m 4307,9693 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7428" />
        <path
           d="m 4391,9566 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7430" />
        <path
           d="m 4601,9247 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7432" />
        <path
           d="m 6707,6067 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7434" />
        <path
           d="m 6833,5875 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7436" />
        <path
           d="m 3794,10123 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7438" />
        <path
           d="m 3738,9936 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7440" />
        <path
           d="m 3613,9513 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7442" />
        <path
           d="m 3525,9215 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7444" />
        <path
           d="m 3469,9028 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7446" />
        <path
           d="m 3943,11617 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7448" />
        <path
           d="m 3855,11319 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7450" />
        <path
           d="m 3800,11132 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7452" />
        <path
           d="m 3674,10709 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7454" />
        <path
           d="m 3586,10411 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7456" />
        <path
           d="m 3531,10224 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7458" />
        <path
           d="m 3406,9801 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7460" />
        <path
           d="m 3317,9503 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7462" />
        <path
           d="m 3137,8893 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7464" />
        <path
           d="m 3055,9604 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7466" />
        <path
           d="m 3736,11905 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7468" />
        <path
           d="m 3648,11607 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7470" />
        <path
           d="m 3592,11420 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7472" />
        <path
           d="m 3467,10997 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7474" />
        <path
           d="m 3379,10699 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7476" />
        <path
           d="m 3323,10512 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7478" />
        <path
           d="m 3198,10089 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7480" />
        <path
           d="m 3110,9791 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7482" />
        <path
           d="m 3529,12193 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7484" />
        <path
           d="m 3440,11895 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7486" />
        <path
           d="m 3385,11708 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7488" />
        <path
           d="m 3260,11285 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7490" />
        <path
           d="m 3171,10987 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7492" />
        <path
           d="m 3116,10800 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7494" />
        <path
           d="m 2991,10378 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7496" />
        <path
           d="m 2903,10080 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7498" />
        <path
           d="m 2847,9893 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7500" />
        <path
           d="m 3321,12481 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7502" />
        <path
           d="m 3233,12183 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7504" />
        <path
           d="m 3178,11996 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7506" />
        <path
           d="m 3052,11574 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7508" />
        <path
           d="m 2964,11276 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7510" />
        <path
           d="m 2909,11089 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7512" />
        <path
           d="m 2783,10666 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7514" />
        <path
           d="m 2695,10368 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7516" />
        <path
           d="m 2640,10181 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7518" />
        <path
           d="m 2576,10954 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7520" />
        <path
           d="m 3114,12770 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7522" />
        <path
           d="m 3026,12472 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7524" />
        <path
           d="m 2970,12285 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7526" />
        <path
           d="m 2845,11862 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7528" />
        <path
           d="m 2757,11564 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7530" />
        <path
           d="m 2701,11377 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7532" />
        <path
           d="m 2488,10656 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7534" />
        <path
           d="m 2432,10469 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7536" />
        <path
           d="m 3032,13481 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7538" />
        <path
           d="m 2906,13058 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7540" />
        <path
           d="m 2818,12760 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7542" />
        <path
           d="m 2763,12573 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7544" />
        <path
           d="m 2638,12150 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7546" />
        <path
           d="m 2549,11852 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7548" />
        <path
           d="m 2494,11665 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7550" />
        <path
           d="m 2369,11242 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7552" />
        <path
           d="m 2280,10944 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7554" />
        <path
           d="m 2225,10757 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7556" />
        <path
           d="m 2824,13769 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7558" />
        <path
           d="m 2699,13346 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7560" />
        <path
           d="m 2611,13048 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7562" />
        <path
           d="m 2555,12861 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7564" />
        <path
           d="m 2430,12438 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7566" />
        <path
           d="m 2342,12140 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7568" />
        <path
           d="m 2287,11953 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7570" />
        <path
           d="m 2161,11530 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7572" />
        <path
           d="m 2073,11232 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7574" />
        <path
           d="m 2018,11045 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7576" />
        <path
           d="m 2492,13634 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7578" />
        <path
           d="m 2403,13336 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7580" />
        <path
           d="m 2348,13149 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7582" />
        <path
           d="m 2223,12726 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7584" />
        <path
           d="m 2135,12428 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7586" />
        <path
           d="m 2079,12241 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7588" />
        <path
           d="m 1954,11818 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7590" />
        <path
           d="m 1866,11520 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7592" />
        <path
           d="m 2196,13624 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7594" />
        <path
           d="m 2141,13437 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7596" />
        <path
           d="m 2015,13014 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7598" />
        <path
           d="m 1927,12716 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7600" />
        <path
           d="m 1872,12530 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7602" />
        <path
           d="m 1746,12107 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7604" />
        <path
           d="m 1658,11809 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7606" />
        <path
           d="m 2202,14633 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7608" />
        <path
           d="m 1989,13913 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7610" />
        <path
           d="m 1933,13726 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7612" />
        <path
           d="m 1808,13303 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7614" />
        <path
           d="m 1720,13005 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7616" />
        <path
           d="m 1664,12818 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7618" />
        <path
           d="m 1539,12395 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7620" />
        <path
           d="m 1451,12097 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7622" />
        <path
           d="m 1870,14499 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7624" />
        <path
           d="m 1781,14201 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7626" />
        <path
           d="m 1726,14014 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7628" />
        <path
           d="m 1601,13591 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7630" />
        <path
           d="m 1512,13293 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7632" />
        <path
           d="m 1457,13106 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7634" />
        <path
           d="m 1332,12683 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7636" />
        <path
           d="m 1519,14302 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7638" />
        <path
           d="m 1393,13879 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7640" />
        <path
           d="m 1305,13581 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7642" />
        <path
           d="m 1250,13394 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7644" />
        <path
           d="m 1124,12971 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7646" />
        <path
           d="m 1098,13869 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7648" />
        <path
           d="m 1042,13682 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7650" />
        <path
           d="m 917,13259 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7652" />
        <path
           d="m 835,13970 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7654" />
        <path
           d="m 710,13548 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7656" />
        <path
           d="m 7178,5589 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7658" />
        <path
           d="m 7050,5883 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7660" />
        <path
           d="m 6851,5559 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7662" />
        <path
           d="m 6723,5853 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7664" />
        <path
           d="m 6595,6147 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7666" />
        <path
           d="m 6542,5682 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7668" />
        <path
           d="m 6525,5533 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7670" />
        <path
           d="m 6414,5976 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7672" />
        <path
           d="m 6397,5827 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7674" />
        <path
           d="m 6198,5504 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7676" />
        <path
           d="m 6070,5797 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7678" />
        <path
           d="m 6017,5332 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7680" />
        <path
           d="m 6012,6708 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7682" />
        <path
           d="m 5942,6091 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7684" />
        <path
           d="m 5889,5626 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7686" />
        <path
           d="m 5872,5477 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7688" />
        <path
           d="m 5884,7002 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7690" />
        <path
           d="m 5813,6385 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7692" />
        <path
           d="m 5760,5920 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7694" />
        <path
           d="m 5743,5771 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7696" />
        <path
           d="m 5825,7910 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7698" />
        <path
           d="m 5755,7296 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7700" />
        <path
           d="m 5685,6679 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7702" />
        <path
           d="m 5632,6214 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7704" />
        <path
           d="m 5615,6065 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7706" />
        <path
           d="m 5545,5448 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7708" />
        <path
           d="m 5697,8204 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7710" />
        <path
           d="m 5644,7739 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7712" />
        <path
           d="m 5627,7590 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7714" />
        <path
           d="m 5557,6973 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7716" />
        <path
           d="m 5504,6508 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7718" />
        <path
           d="m 5487,6359 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7720" />
        <path
           d="m 5417,5742 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7722" />
        <path
           d="m 5569,8498 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7724" />
        <path
           d="m 5516,8033 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7726" />
        <path
           d="m 5499,7884 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7728" />
        <path
           d="m 5429,7267 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7730" />
        <path
           d="m 5376,6802 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7732" />
        <path
           d="m 5359,6653 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7734" />
        <path
           d="m 5288,6035 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7736" />
        <path
           d="m 5235,5570 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7738" />
        <path
           d="m 5441,8791 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7740" />
        <path
           d="m 5388,8326 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7742" />
        <path
           d="m 5371,8177 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7744" />
        <path
           d="m 5300,7560 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7746" />
        <path
           d="m 5247,7095 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7748" />
        <path
           d="m 5230,6946 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7750" />
        <path
           d="m 5160,6329 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7752" />
        <path
           d="m 5107,5864 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7754" />
        <path
           d="m 5090,5715 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7756" />
        <path
           d="m 5172,7854 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7758" />
        <path
           d="m 5119,7389 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7760" />
        <path
           d="m 5102,7240 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7762" />
        <path
           d="m 5032,6623 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7764" />
        <path
           d="m 4979,6158 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7766" />
        <path
           d="m 4962,6009 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7768" />
        <path
           d="m 5312,9085 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7770" />
        <path
           d="m 5044,8148 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7772" />
        <path
           d="m 4991,7683 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7774" />
        <path
           d="m 4974,7534 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7776" />
        <path
           d="m 4904,6917 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7778" />
        <path
           d="m 4851,6452 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7780" />
        <path
           d="m 4834,6303 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7782" />
        <path
           d="m 4916,8442 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7784" />
        <path
           d="m 4863,7977 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7786" />
        <path
           d="m 4846,7828 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7788" />
        <path
           d="m 4775,7211 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7790" />
        <path
           d="m 4722,6746 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7792" />
        <path
           d="m 4705,6597 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7794" />
        <path
           d="m 4635,5980 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7796" />
        <path
           d="m 4787,8736 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7798" />
        <path
           d="m 4734,8271 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7800" />
        <path
           d="m 4717,8122 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7802" />
        <path
           d="m 4647,7505 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7804" />
        <path
           d="m 4594,7040 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7806" />
        <path
           d="m 4577,6891 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7808" />
        <path
           d="m 4507,6274 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7810" />
        <path
           d="m 4659,9029 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7812" />
        <path
           d="m 4606,8564 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7814" />
        <path
           d="m 4589,8415 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7816" />
        <path
           d="m 4519,7798 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7818" />
        <path
           d="m 4466,7333 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7820" />
        <path
           d="m 4449,7184 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7822" />
        <path
           d="m 4379,6567 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7824" />
        <path
           d="m 4531,9323 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7826" />
        <path
           d="m 4478,8858 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7828" />
        <path
           d="m 4461,8709 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7830" />
        <path
           d="m 4391,8092 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7832" />
        <path
           d="m 4338,7627 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7834" />
        <path
           d="m 4321,7478 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7836" />
        <path
           d="m 4618,10089 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7838" />
        <path
           d="m 4601,9940 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7840" />
        <path
           d="m 4250,6861 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7842" />
        <path
           d="m 4490,10383 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7844" />
        <path
           d="m 4473,10234 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7846" />
        <path
           d="m 4403,9617 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7848" />
        <path
           d="m 4350,9152 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7850" />
        <path
           d="m 4333,9003 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7852" />
        <path
           d="m 4262,8386 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7854" />
        <path
           d="m 4209,7921 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7856" />
        <path
           d="m 4192,7772 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7858" />
        <path
           d="m 4122,7155 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7860" />
        <path
           d="m 4345,10528 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7862" />
        <path
           d="m 4274,9911 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7864" />
        <path
           d="m 4221,9446 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7866" />
        <path
           d="m 4204,9297 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7868" />
        <path
           d="m 4134,8680 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7870" />
        <path
           d="m 4081,8215 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7872" />
        <path
           d="m 4064,8066 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7874" />
        <path
           d="m 3994,7449 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7876" />
        <path
           d="m 4146,10205 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7878" />
        <path
           d="m 4093,9740 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7880" />
        <path
           d="m 4076,9591 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7882" />
        <path
           d="m 4006,8974 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7884" />
        <path
           d="m 3953,8509 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7886" />
        <path
           d="m 3936,8360 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7888" />
        <path
           d="m 4233,10971 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7890" />
        <path
           d="m 4216,10822 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7892" />
        <path
           d="m 4018,10499 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7894" />
        <path
           d="m 3965,10034 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7896" />
        <path
           d="m 3948,9885 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7898" />
        <path
           d="m 3878,9267 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7900" />
        <path
           d="m 3825,8802 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7902" />
        <path
           d="m 3808,8653 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7904" />
        <path
           d="m 4105,11265 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7906" />
        <path
           d="m 4088,11116 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7908" />
        <path
           d="m 3977,11558 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7910" />
        <path
           d="m 3960,11409 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7912" />
        <path
           d="m 3890,10792 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7914" />
        <path
           d="m 3837,10327 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7916" />
        <path
           d="m 3820,10178 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7918" />
        <path
           d="m 3749,9561 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7920" />
        <path
           d="m 3696,9096 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7922" />
        <path
           d="m 3679,8947 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7924" />
        <path
           d="m 3481,8624 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7926" />
        <path
           d="m 3849,11852 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7928" />
        <path
           d="m 3832,11703 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7930" />
        <path
           d="m 3761,11086 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7932" />
        <path
           d="m 3708,10621 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7934" />
        <path
           d="m 3691,10472 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7936" />
        <path
           d="m 3621,9855 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7938" />
        <path
           d="m 3568,9390 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7940" />
        <path
           d="m 3551,9241 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7942" />
        <path
           d="m 3353,8918 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7944" />
        <path
           d="m 3720,12146 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7946" />
        <path
           d="m 3703,11997 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7948" />
        <path
           d="m 6904,5800 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7950" />
        <path
           d="m 6849,5613 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7952" />
        <path
           d="m 6697,6088 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7954" />
        <path
           d="m 6642,5901 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7956" />
        <path
           d="m 6516,5479 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7958" />
        <path
           d="m 6309,5767 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7960" />
        <path
           d="m 6221,5469 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7962" />
        <path
           d="m 6370,6963 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7964" />
        <path
           d="m 6102,6055 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7966" />
        <path
           d="m 6013,5757 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7968" />
        <path
           d="m 5958,5570 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7970" />
        <path
           d="m 6163,7251 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7972" />
        <path
           d="m 6019,6766 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7974" />
        <path
           d="m 5894,6343 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7976" />
        <path
           d="m 5806,6045 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7978" />
        <path
           d="m 5750,5858 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7980" />
        <path
           d="m 5625,5435 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7982" />
        <path
           d="m 5812,7054 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7984" />
        <path
           d="m 5687,6631 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7986" />
        <path
           d="m 5598,6333 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7988" />
        <path
           d="m 5543,6146 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7990" />
        <path
           d="m 5418,5723 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7992" />
        <path
           d="m 5330,5425 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7994" />
        <path
           d="m 5748,7827 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7996" />
        <path
           d="m 5660,7529 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path7998" />
        <path
           d="m 5605,7342 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8000" />
        <path
           d="m 5479,6919 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8002" />
        <path
           d="m 5391,6621 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8004" />
        <path
           d="m 5336,6434 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8006" />
        <path
           d="m 5210,6012 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8008" />
        <path
           d="m 5122,5714 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8010" />
        <path
           d="m 5067,5527 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8012" />
        <path
           d="m 5541,8115 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8014" />
        <path
           d="m 5453,7817 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8016" />
        <path
           d="m 5397,7630 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8018" />
        <path
           d="m 5272,7208 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8020" />
        <path
           d="m 5184,6910 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8022" />
        <path
           d="m 5128,6723 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8024" />
        <path
           d="m 5003,6300 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8026" />
        <path
           d="m 4859,5815 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8028" />
        <path
           d="m 5245,8106 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8030" />
        <path
           d="m 5190,7919 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8032" />
        <path
           d="m 5065,7496 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8034" />
        <path
           d="m 4976,7198 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8036" />
        <path
           d="m 4921,7011 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8038" />
        <path
           d="m 4796,6588 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8040" />
        <path
           d="m 5459,8827 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8042" />
        <path
           d="m 4652,6103 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8044" />
        <path
           d="m 5038,8394 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8046" />
        <path
           d="m 4982,8207 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8048" />
        <path
           d="m 4857,7784 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8050" />
        <path
           d="m 4769,7486 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8052" />
        <path
           d="m 4714,7299 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8054" />
        <path
           d="m 4588,6876 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8056" />
        <path
           d="m 5251,9115 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8058" />
        <path
           d="m 4445,6391 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8060" />
        <path
           d="m 4830,8682 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8062" />
        <path
           d="m 4775,8495 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8064" />
        <path
           d="m 4650,8072 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8066" />
        <path
           d="m 4562,7774 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8068" />
        <path
           d="m 4506,7587 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8070" />
        <path
           d="m 4293,6866 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8072" />
        <path
           d="m 4623,8970 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8074" />
        <path
           d="m 4568,8783 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8076" />
        <path
           d="m 4442,8360 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8078" />
        <path
           d="m 4354,8062 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8080" />
        <path
           d="m 4299,7875 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8082" />
        <path
           d="m 4174,7453 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8084" />
        <path
           d="m 4085,7155 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8086" />
        <path
           d="m 4416,9258 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8088" />
        <path
           d="m 4360,9071 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8090" />
        <path
           d="m 4235,8649 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8092" />
        <path
           d="m 4147,8351 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8094" />
        <path
           d="m 4091,8164 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8096" />
        <path
           d="m 4685,10166 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8098" />
        <path
           d="m 4629,9979 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8100" />
        <path
           d="m 3966,7741 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8102" />
        <path
           d="m 3878,7443 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8104" />
        <path
           d="m 4477,10454 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8106" />
        <path
           d="m 4422,10267 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8108" />
        <path
           d="m 4297,9845 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8110" />
        <path
           d="m 4208,9547 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8112" />
        <path
           d="m 4153,9360 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8114" />
        <path
           d="m 4028,8937 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8116" />
        <path
           d="m 3939,8639 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8118" />
        <path
           d="m 3884,8452 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8120" />
        <path
           d="m 4089,10133 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8122" />
        <path
           d="m 4001,9835 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8124" />
        <path
           d="m 3946,9648 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8126" />
        <path
           d="m 3820,9225 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8128" />
        <path
           d="m 3732,8927 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8130" />
        <path
           d="m 3677,8740 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8132" />
        <path
           d="m 3344,8605 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8134" />
        <path
           d="m 4151,11329 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8136" />
        <path
           d="m 4062,11031 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8138" />
        <path
           d="m 4007,10844 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8140" />
        <path
           d="m 3882,10421 v 0"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:0.74902"
           id="path8142" />
        <path
           d="m 6108,6698 265,140 -418,797 -266,-140 419,-797"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8144" />
        <path
           d="m 4826,9137 266,140 418,-797 -265,-140 -419,797"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8146" />
        <path
           d="m 6615,6503 74,39 -58,112 -75,-39 59,-112"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8148" />
        <path
           d="m 4887,9512.5 c 0,30.6514 -24.8481,55.5 -55.5,55.5 -30.6519,0 -55.5,-24.8486 -55.5,-55.5 0,-30.6514 24.8481,-55.5 55.5,-55.5 30.6519,0 55.5,24.8486 55.5,55.5"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8150" />
        <path
           d="m 4828,10848 299,157 -105,199 -298,-157 104,-199"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8152" />
        <path
           d="m 4142,10479 299,157 -105,199 -299,-157 105,-199"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8154" />
        <path
           d="m 4145,10490 285,150 -97,185 -285,-150 97,-185"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8156" />
        <path
           d="m 4363,10709 -1,5 -1,5 -2,4 -3,4 -4,3 -4,2 -5,2 -4,1 -5,-1 -5,-1 -4,-2 -4,-3 -4,-3 -2,-4 -2,-5 -1,-4 v -5 l 1,-5 2,-5 2,-4 4,-3 4,-3 4,-2 5,-1 h 5 4 l 5,2 4,2 4,3 3,4 2,5 1,4 1,5"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8158" />
        <path
           d="m 4166,10606 v 4 l -2,5 -2,4 -3,4 -4,3 -4,3 -4,1 -5,1 h -5 l -5,-1 -4,-2 -4,-3 -3,-4 -3,-4 -2,-4 -1,-5 v -5 l 1,-5 2,-4 3,-4 3,-4 4,-2 4,-2 5,-2 h 5 l 5,1 4,1 4,3 4,3 3,4 2,4 2,5 v 5"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8160" />
        <path
           d="m 5239,5280 99,5 36,-30 -30,70 -93,-1 54,65 39,6 -46,21 -64,-72 -53,87 -80,6 68,-22 42,-98 -113,-53 -29,26 25,-57 110,31 22,-93 -26,-13 61,13 -22,109"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8162" />
        <path
           d="m 5112,5254 123,50"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8164" />
        <path
           d="m 5178,5419 58,-115"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8166" />
        <path
           d="m 5232,5311 64,88"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8168" />
        <path
           d="m 5231,5304 100,2"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8170" />
        <path
           d="m 5231,5302 -6,-25 15,-94"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8172" />
        <path
           d="m 5348,5300.5 c 0,64.8935 -52.6065,117.5 -117.5,117.5 -64.8936,0 -117.5,-52.6065 -117.5,-117.5 0,-64.8936 52.6064,-117.5 117.5,-117.5 64.8935,0 117.5,52.6064 117.5,117.5"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8174" />
        <path
           d="m 5359,5300.5 c 0,70.9687 -57.5313,128.5 -128.5,128.5 -70.9688,0 -128.5,-57.5313 -128.5,-128.5 0,-70.9688 57.5312,-128.5 128.5,-128.5 70.9687,0 128.5,57.5312 128.5,128.5"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8176" />
        <path
           d="m 3350,8686 99,5 37,-30 -30,70 -94,-1 55,65 39,6 -47,21 -64,-72 -52,86 -81,7 68,-23 43,-97 -114,-53 -28,26 24,-57 111,31 21,-93 -25,-13 60,12 -22,110"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8178" />
        <path
           d="m 3224,8660 122,50"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8180" />
        <path
           d="m 3290,8825 57,-115"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8182" />
        <path
           d="m 3344,8717 64,87"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8184" />
        <path
           d="m 3343,8710 99,1"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8186" />
        <path
           d="m 3342,8708 -6,-25 16,-94"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8188" />
        <path
           d="m 3460,8705.5 c 0,64.8936 -52.6064,117.5 -117.5,117.5 -64.8936,0 -117.5,-52.6064 -117.5,-117.5 0,-64.8935 52.6064,-117.5 117.5,-117.5 64.8936,0 117.5,52.6065 117.5,117.5"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8190" />
        <path
           d="m 3471,8705.5 c 0,70.9688 -57.5315,128.5 -128.5,128.5 -70.9685,0 -128.5,-57.5312 -128.5,-128.5 0,-70.9687 57.5315,-128.5 128.5,-128.5 70.9685,0 128.5,57.5313 128.5,128.5"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8192" />
        <path
           d="m 912,12986 967,508"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8194" />
        <path
           d="m 2045,13581 166,88"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8196" />
        <path
           d="m 2377,13756 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8198" />
        <path
           d="m 2709,13930 830,436"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8200" />
        <path
           d="m 3705,14453 166,88"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8202" />
        <path
           d="m 4037,14628 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8204" />
        <path
           d="m 4369,14802 968,509"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8206" />
        <path
           d="m 587,13680 952,500"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8208" />
        <path
           d="m 1705,14267 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8210" />
        <path
           d="m 2037,14441 166,88"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8212" />
        <path
           d="m 2369,14616 830,436"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8214" />
        <path
           d="m 3365,15139 166,87"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8216" />
        <path
           d="m 3697,15313 166,88"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8218" />
        <path
           d="m 4029,15488 952,500"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8220" />
        <path
           d="m 593,16380 181,48"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8222" />
        <path
           d="m 955,16477 705,188 608,320"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8224" />
        <path
           d="m 2434,17072 166,88"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8226" />
        <path
           d="m 2766,17247 166,87"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8228" />
        <path
           d="m 3098,17421 830,436"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8230" />
        <path
           d="m 4094,17944 166,88"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8232" />
        <path
           d="m 4426,18119 166,87"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8234" />
        <path
           d="m 4758,18293 830,436"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8236" />
        <path
           d="m 5754,18816 166,87"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8238" />
        <path
           d="m 10263,17356 605,343"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8240" />
        <path
           d="m 11031,17792 164,92"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8242" />
        <path
           d="m 11358,17977 163,92"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8244" />
        <path
           d="m 11684,18162 519,294"
           style="fill:none;stroke:#00a5dd;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8246" />
        <path
           d="m 3310,9421.5 c 0,104.1055 -84.3943,188.5 -188.5,188.5 -104.1057,0 -188.5,-84.3945 -188.5,-188.5 0,-104.1055 84.3943,-188.5 188.5,-188.5 104.1057,0 188.5,84.3945 188.5,188.5"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8248" />
        <path
           d="m 3131,9129 106,-202 208,109 -106,202 -208,-109"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8250" />
        <path
           d="m 2886,9595 -106,202 208,109 106,-202 -208,-109"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8252" />
        <path
           d="m 3441,8409 199,105 384,-730 -200,-105 -383,730"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8254" />
        <path
           d="m 4120,7116 266,139 122,-232 -266,-140 -122,233"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8256" />
        <path
           d="m 4772,5875 199,105 -384,730 -199,-104 384,-731"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8258" />
        <path
           d="m 1474,13281 93,-176"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8260" />
        <path
           d="m 1610,13022 88,-166"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8262" />
        <path
           d="m 1741,12773 87,-166"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8264" />
        <path
           d="m 1872,12524 87,-166"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8266" />
        <path
           d="m 2003,12275 87,-166"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8268" />
        <path
           d="m 2134,12026 87,-166"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8270" />
        <path
           d="m 2264,11777 88,-166"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8272" />
        <path
           d="m 2395,11528 87,-166"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8274" />
        <path
           d="m 2526,11279 93,-176 -44,-139"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8276" />
        <path
           d="m 2547,10874 -43,-139 -103,-54"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8278" />
        <path
           d="m 2318,10637 -104,-54"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8280" />
        <path
           d="m 4285,7418.5 c 0,20.7104 -16.7896,37.5 -37.5,37.5 -20.7105,0 -37.5,-16.7896 -37.5,-37.5 0,-20.7105 16.7895,-37.5 37.5,-37.5 20.7104,0 37.5,16.7895 37.5,37.5"
           style="fill:none;stroke:#000000;stroke-width:24;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8282" />
        <path
           d="m 4525,8191.5 c 0,20.7109 -16.7896,37.5 -37.5,37.5 -20.7105,0 -37.5,-16.7891 -37.5,-37.5 0,-20.7105 16.7895,-37.5 37.5,-37.5 20.7104,0 37.5,16.7895 37.5,37.5"
           style="fill:none;stroke:#000000;stroke-width:24;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8284" />
        <path
           d="m 2542,10735.5 c 0,20.711 -16.7893,37.5 -37.5,37.5 -20.7107,0 -37.5,-16.789 -37.5,-37.5 0,-20.711 16.7893,-37.5 37.5,-37.5 20.7107,0 37.5,16.789 37.5,37.5"
           style="fill:none;stroke:#808080;stroke-width:24;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8286" />
        <path
           d="m 2657,11103.5 c 0,20.711 -16.7893,37.5 -37.5,37.5 -20.7107,0 -37.5,-16.789 -37.5,-37.5 0,-20.711 16.7893,-37.5 37.5,-37.5 20.7107,0 37.5,16.789 37.5,37.5"
           style="fill:none;stroke:#808080;stroke-width:24;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8288" />
        <path
           d="M 1740,13421 4487,8191 4247,7418 3957,7265"
           style="fill:none;stroke:#000000;stroke-width:24;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8290" />
        <path
           d="m 518,13812 4586,-8731 2129,463 -421,801 -531,-279 -279,531 531,279 -1318,2511 -532,-279 -279,531 532,279 -2559,4871 -1859,-977"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8292" />
        <path
           d="m 9275,14040 361,190"
           style="fill:none;stroke:#ff0000;stroke-width:14;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8294" />
        <path
           d="m 2201,13833 532,279 -279,531 -532,-279 279,-531"
           style="fill:none;stroke:#0000ff;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8296" />
        <path
           d="m 1735.57,14287.734 c -89.2593,-44.309 -135.9946,-144.472 -112.6067,-241.341 23.3877,-96.869 110.6771,-164.674 210.3204,-163.374"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8298" />
        <path
           d="m 1833.5127,13882.93 c -52.99,-96.671 -27.5771,-217.54 59.8555,-284.688 87.4326,-67.147 210.7668,-60.513 290.4922,15.625"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8300" />
        <path
           d="m 2182.7813,13614.145 c 25.8388,-98.073 119.3613,-162.629 220.2236,-152.017 100.862,10.613 178.8992,93.223 183.759,194.524"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8302" />
        <path
           d="m 2587.3071,13656.72 c 68.1531,-55.812 167.1197,-52.454 231.333,7.848 64.2137,60.303 73.7754,158.864 22.3509,230.385"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8304" />
        <path
           d="m 2841.5022,13896.006 c 128.9272,-17.699 255.9082,43.58 322.2722,155.522 66.3643,111.944 59.1895,252.755 -18.209,357.373 -77.3987,104.619 -209.9506,152.673 -336.4111,121.961"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8306" />
        <path
           d="m 2809.0666,14530.369 c 37.9612,55.422 42.4068,127.218 11.5723,186.9 -30.8342,59.681 -91.9626,97.598 -159.1296,98.707"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8308" />
        <path
           d="m 2661.8945,14815.776 c -44.9751,157.115 -203.1001,253.325 -363.3068,221.05 -160.2068,-32.274 -268.7458,-182.205 -249.3785,-344.478"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8310" />
        <path
           d="m 2049.4202,14692.449 c -112.2458,77.644 -265.6361,53.792 -349.0054,-54.269 -83.3694,-108.062 -67.5171,-262.484 36.0684,-351.353"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8312" />
        <path
           d="m 2405,14236.5 c 0,30.651 -24.8481,55.5 -55.5,55.5 -30.6519,0 -55.5,-24.849 -55.5,-55.5 0,-30.651 24.8481,-55.5 55.5,-55.5 30.6519,0 55.5,24.849 55.5,55.5"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8314" />
        <path
           d="m 2454,14643 -532,-279 279,-531 532,279"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8316" />
        <path
           d="m 1512,13281.5 c 0,20.711 -16.7893,37.5 -37.5,37.5 -20.7107,0 -37.5,-16.789 -37.5,-37.5 0,-20.711 16.7893,-37.5 37.5,-37.5 20.7107,0 37.5,16.789 37.5,37.5"
           style="fill:none;stroke:#808080;stroke-width:24;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8318" />
        <path
           d="m 1157,13959.5 c 0,20.711 -16.7893,37.5 -37.5,37.5 -20.7107,0 -37.5,-16.789 -37.5,-37.5 0,-20.711 16.7893,-37.5 37.5,-37.5 20.7107,0 37.5,16.789 37.5,37.5"
           style="fill:none;stroke:#808080;stroke-width:24;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8320" />
      </g>
    </g>
    <g
       id="g8322">
      <g
         id="g8324"
         clip-path="url(#clipPath8328)">
        <g
           id="g8330">
          <path
             d="m 12029,18180 h -600 l 600,-90 z m -600,0 600,-90 h -600 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8332" />
        </g>
        <g
           id="g8334">
          <path
             d="m 10829,18180 h -300 l 300,-90 z m -300,0 300,-90 h -300 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8336" />
        </g>
        <g
           id="g8338">
          <path
             d="m 10229,18180 h -300 l 300,-90 z m -300,0 300,-90 h -300 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8340" />
        </g>
        <g
           id="g8342">
          <path
             d="m 11429,18090 h -600 l 600,-90 z m -600,0 600,-90 h -600 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8344" />
        </g>
        <g
           id="g8346">
          <path
             d="m 10529,18090 h -300 l 300,-90 z m -300,0 300,-90 h -300 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8348" />
        </g>
        <g
           id="g8350">
          <path
             d="m 9929,18090 h -300 l 300,-90 z m -300,0 300,-90 h -300 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8352" />
        </g>
        <path
           d="m 10249,17838 -11,14 -15,7 h -21 l -15,-7 -10,-14 v -13 l 5,-14 5,-7 10,-7 31,-14 10,-6 6,-7 5,-14 v -21 l -11,-13 -15,-7 h -21 l -15,7 -10,13"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8354" />
        <path
           d="m 10357,17825 -5,13 -11,14 -10,7 h -21 l -10,-7 -10,-14 -5,-13 -5,-21 v -34 l 5,-21 5,-14 10,-13 10,-7 h 21 l 10,7 11,13 5,14"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8356" />
        <path
           d="m 10388,17715 41,144 41,-144"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8358" />
        <path
           d="m 10403,17763 h 51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8360" />
        <path
           d="m 10501,17859 v -144 h 61"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8362" />
        <path
           d="m 10588,17715 v 144 h 67"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8364" />
        <path
           d="m 10588,17790 h 41"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8366" />
        <path
           d="m 10588,17715 h 67"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8368" />
        <path
           d="m 10691,17811 -5,-7 5,-7 5,7 -5,7"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8370" />
        <path
           d="m 10691,17729 -5,-7 5,-7 5,7 -5,7"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8372" />
        <path
           d="m 10861,17831 10,7 15,21 v -144"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8374" />
        <path
           d="m 10953,17879 -5,-6 -5,6 5,7 5,-7 v -13 l -5,-14 -5,-7"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8376" />
        <path
           d="m 10984,17879 -5,-6 -5,6 5,7 5,-7 v -13 l -5,-14 -5,-7"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8378" />
        <path
           d="m 11118,17797 h 92"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8380" />
        <path
           d="m 11118,17756 h 92"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8382" />
        <path
           d="m 11375,17859 -15,-7 -6,-14 v -13 l 6,-14 10,-7 20,-7 16,-7 10,-13 5,-14 v -21 l -5,-13 -5,-7 -15,-7 h -21 l -15,7 -6,7 -5,13 v 21 l 5,14 11,13 15,7 21,7 10,7 5,14 v 13 l -5,14 -15,7 h -21"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8384" />
        <path
           d="m 11462,17879 -5,-6 -5,6 5,7 5,-7 v -13 l -5,-14 -5,-7"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8386" />
        <path
           d="m 10820,18765 v -508"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8388" />
        <path
           d="m 10759,18646 61,119 57,-119"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8390" />
        <path
           d="m 10755,18360 v 134 l 140,-139 v 139"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8392" />
        <path
           d="m 9629,18000 v 180 h 2400 v -180 H 9629"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8394" />
        <path
           d="m 10829,18180 v -180"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8396" />
        <path
           d="m 10229,18180 v -180"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8398" />
        <path
           d="m 9929,18180 v -180"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8400" />
        <path
           d="m 10529,18180 v -180"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8402" />
        <path
           d="m 11429,18180 v -180"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8404" />
        <path
           d="m 9629,18090 h 2400"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8406" />
        <path
           d="M 8,5 H 12649 V 19378 H 8 V 5"
           style="fill:none;stroke:#767676;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path8408" />
        <g
           id="g8410">
          <path
             d="m 459,18928 -12,12 12,-18469 z m -12,12 L 459,471 447,459 Z M 459,471 447,459 12198,471 Z m -12,-12 11751,12 12,-12 z m 11751,12 12,-12 -12,18469 z m 12,-12 -12,18469 12,12 z m -12,18469 12,12 -11751,-12 z m 12,12 -11751,-12 -12,12 z"
             style="fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:#0000ff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8412" />
        </g>
        <g
           id="g8414">
          <path
             d="M 811,1513 H 703 l 108,-8 z m -108,0 108,-8 H 703 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8416" />
        </g>
        <g
           id="g8418">
          <path
             d="m 725,1505 v 0 h -22 z m 0,0 h -22 28 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8420" />
        </g>
        <g
           id="g8422">
          <path
             d="m 811,1505 h -27 l 27,-1 z m -27,0 27,-1 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8424" />
        </g>
        <g
           id="g8426">
          <path
             d="m 725,1505 h -22 l 17,-1 z m -22,0 17,-1 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8428" />
        </g>
        <g
           id="g8430">
          <path
             d="m 811,1504 h -21 l 21,-1 z m -21,0 21,-1 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8432" />
        </g>
        <g
           id="g8434">
          <path
             d="m 720,1504 h -18 l 15,-1 z m -18,0 15,-1 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8436" />
        </g>
        <g
           id="g8438">
          <path
             d="m 811,1503 h -16 l 16,-2 z m -16,0 16,-2 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8440" />
        </g>
        <g
           id="g8442">
          <path
             d="m 717,1503 h -15 l 11,-2 z m -15,0 11,-2 h -11 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8444" />
        </g>
        <g
           id="g8446">
          <path
             d="m 811,1501 h -12 l 12,-2 z m -12,0 12,-2 h -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8448" />
        </g>
        <g
           id="g8450">
          <path
             d="m 713,1501 h -11 l 8,-3 z m -11,0 8,-3 h -8 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8452" />
        </g>
        <g
           id="g8454">
          <path
             d="m 811,1499 h -9 l 10,-4 z m -9,0 10,-4 h -7 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8456" />
        </g>
        <g
           id="g8458">
          <path
             d="m 710,1498 h -8 l 6,-5 z m -8,0 6,-5 h -6 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8460" />
        </g>
        <g
           id="g8462">
          <path
             d="m 812,1495 h -7 l 7,-3 z m -7,0 7,-3 h -6 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8464" />
        </g>
        <g
           id="g8466">
          <path
             d="m 708,1493 h -6 l 4,-5 z m -6,0 4,-5 h -4 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8468" />
        </g>
        <g
           id="g8470">
          <path
             d="m 812,1492 h -6 l 6,-4 z m -6,0 6,-4 h -4 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8472" />
        </g>
        <g
           id="g8474">
          <path
             d="m 812,1488 h -4 l 4,-6 z m -4,0 4,-6 h -4 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8476" />
        </g>
        <g
           id="g8478">
          <path
             d="m 706,1488 h -4 l 3,-6 z m -4,0 3,-6 h -4 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8480" />
        </g>
        <g
           id="g8482">
          <path
             d="m 766,1505 h -19 l 19,-101 z m -19,0 19,-101 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8484" />
        </g>
        <g
           id="g8486">
          <path
             d="m 766,1404 h -19 l 19,-5 z m -19,0 19,-5 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8488" />
        </g>
        <g
           id="g8490">
          <path
             d="m 766,1399 h -19 l 19,-1 z m -19,0 19,-1 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8492" />
        </g>
        <g
           id="g8494">
          <path
             d="m 766,1398 h -19 l 19,-3 z m -19,0 19,-3 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8496" />
        </g>
        <g
           id="g8498">
          <path
             d="m 766,1395 h -19 l 19,-1 z m -19,0 19,-1 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8500" />
        </g>
        <g
           id="g8502">
          <path
             d="m 766,1394 h -20 l 21,-2 z m -20,0 21,-2 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8504" />
        </g>
        <g
           id="g8506">
          <path
             d="m 767,1392 h -21 l 21,-1 z m -21,0 21,-1 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8508" />
        </g>
        <g
           id="g8510">
          <path
             d="m 767,1391 h -22 l 23,-1 z m -22,0 23,-1 h -23 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8512" />
        </g>
        <g
           id="g8514">
          <path
             d="m 768,1390 h -23 l 23,-1 z m -23,0 23,-1 h -24 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8516" />
        </g>
        <g
           id="g8518">
          <path
             d="m 768,1389 h -24 l 29,-3 z m -24,0 29,-3 h -33 z m 29,-3 h -33 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8520" />
        </g>
        <g
           id="g8522">
          <path
             d="m 740,1386 h 33 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8524" />
        </g>
        <g
           id="g8526">
          <path
             d="m 773,1386 h -34 l 41,-1 z m -34,0 41,-1 h -47 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8528" />
        </g>
        <g
           id="g8530">
          <path
             d="m 784,1385 h -56 l 56,-4 z m -56,0 56,-4 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8532" />
        </g>
        <g
           id="g8534">
          <path
             d="m 850,1520 h -5 l 5,-11 z m -5,0 5,-11 h -31 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8536" />
        </g>
        <g
           id="g8538">
          <path
             d="m 850,1509 h -31 l 31,-2 z m -31,0 31,-2 h -31 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8540" />
        </g>
        <g
           id="g8542">
          <path
             d="m 850,1507 h -23 l 23,-1 z m -23,0 23,-1 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8544" />
        </g>
        <g
           id="g8546">
          <path
             d="m 827,1507 h -8 l 5,-1 z m -8,0 5,-1 h -5 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8548" />
        </g>
        <g
           id="g8550">
          <path
             d="m 820,1505 h 1 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8552" />
        </g>
        <g
           id="g8554">
          <path
             d="m 850,1506 h -22 l 22,-1 z m -22,0 22,-1 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8556" />
        </g>
        <g
           id="g8558">
          <path
             d="m 824,1506 h -5 l 2,-1 z m -5,0 2,-1 h -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8560" />
        </g>
        <g
           id="g8562">
          <path
             d="m 850,1505 h -19 l 19,-1 z m -19,0 19,-1 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8564" />
        </g>
        <g
           id="g8566">
          <path
             d="m 850,1504 h -18 l 18,-3 z m -18,0 18,-3 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8568" />
        </g>
        <g
           id="g8570">
          <path
             d="m 850,1501 h -17 l 17,-3 z m -17,0 17,-3 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8572" />
        </g>
        <g
           id="g8574">
          <path
             d="m 850,1498 h -17 l 17,-4 z m -17,0 17,-4 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8576" />
        </g>
        <g
           id="g8578">
          <path
             d="m 850,1494 h -17 l 17,-5 z m -17,0 17,-5 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8580" />
        </g>
        <g
           id="g8582">
          <path
             d="m 850,1489 h -17 l 17,-7 z m -17,0 17,-7 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8584" />
        </g>
        <g
           id="g8586">
          <path
             d="m 878,1473 9,-1 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8588" />
        </g>
        <g
           id="g8590">
          <path
             d="m 887,1472 h -13 l 14,-1 z m -13,0 14,-1 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8592" />
        </g>
        <g
           id="g8594">
          <path
             d="m 888,1471 h -18 l 21,-2 z m -18,0 21,-2 h -25 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8596" />
        </g>
        <g
           id="g8598">
          <path
             d="m 891,1469 h -25 l 28,-1 z m -25,0 28,-1 h -30 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8600" />
        </g>
        <g
           id="g8602">
          <path
             d="m 894,1468 h -30 l 31,-2 z m -30,0 31,-2 h -34 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8604" />
        </g>
        <g
           id="g8606">
          <path
             d="m 895,1466 h -34 l 36,-2 z m -34,0 36,-2 h -37 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8608" />
        </g>
        <g
           id="g8610">
          <path
             d="m 897,1464 h -37 l 38,-3 z m -37,0 38,-3 h -42 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8612" />
        </g>
        <g
           id="g8614">
          <path
             d="m 898,1461 h -27 28 z m -27,0 h 28 -26 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8616" />
        </g>
        <g
           id="g8618">
          <path
             d="m 870,1461 v 0 h -14 z m 0,0 h -14 15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8620" />
        </g>
        <g
           id="g8622">
          <path
             d="m 899,1461 h -26 z m -26,0 h 26 -23 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8624" />
        </g>
        <g
           id="g8626">
          <path
             d="m 899,1461 h -23 l 23,-1 z m -23,0 23,-1 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8628" />
        </g>
        <g
           id="g8630">
          <path
             d="m 870,1461 h -14 l 9,-1 z m -14,0 9,-1 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8632" />
        </g>
        <g
           id="g8634">
          <path
             d="m 899,1460 h -21 l 22,-2 z m -21,0 22,-2 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8636" />
        </g>
        <g
           id="g8638">
          <path
             d="m 865,1460 h -10 l 3,-4 z m -10,0 3,-4 h -7 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8640" />
        </g>
        <g
           id="g8642">
          <path
             d="m 850,1482 h -16 l 16,-26 z m -16,0 16,-26 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8644" />
        </g>
        <g
           id="g8646">
          <path
             d="m 858,1456 h -7 l 5,-2 z m -7,0 5,-2 h -6 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8648" />
        </g>
        <g
           id="g8650">
          <path
             d="m 850,1456 h -16 l 16,-2 z m -16,0 16,-2 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8652" />
        </g>
        <g
           id="g8654">
          <path
             d="m 900,1458 h -19 l 20,-4 z m -19,0 20,-4 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8656" />
        </g>
        <g
           id="g8658">
          <path
             d="m 856,1454 h -22 l 20,-1 z m -22,0 20,-1 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8660" />
        </g>
        <g
           id="g8662">
          <path
             d="m 901,1454 h -17 l 17,-3 z m -17,0 17,-3 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8664" />
        </g>
        <g
           id="g8666">
          <path
             d="m 901,1451 h -16 l 17,-2 z m -16,0 17,-2 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8668" />
        </g>
        <g
           id="g8670">
          <path
             d="m 854,1453 h -20 l 16,-5 z m -20,0 16,-5 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8672" />
        </g>
        <g
           id="g8674">
          <path
             d="m 902,1449 h -17 l 17,-2 z m -17,0 17,-2 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8676" />
        </g>
        <g
           id="g8678">
          <path
             d="m 902,1447 h -16 l 16,-5 z m -16,0 16,-5 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8680" />
        </g>
        <g
           id="g8682">
          <path
             d="m 902,1442 h -16 l 16,-1 z m -16,0 16,-1 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8684" />
        </g>
        <g
           id="g8686">
          <path
             d="m 902,1441 h -16 l 16,-8 z m -16,0 16,-8 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8688" />
        </g>
        <g
           id="g8690">
          <path
             d="m 903,1433 v 0 h -17 z m 0,0 h -17 16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8692" />
        </g>
        <g
           id="g8694">
          <path
             d="m 903,1433 h -17 l 17,-32 z m -17,0 17,-32 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8696" />
        </g>
        <g
           id="g8698">
          <path
             d="m 850,1448 h -16 l 16,-47 z m -16,0 16,-47 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8700" />
        </g>
        <g
           id="g8702">
          <path
             d="m 903,1401 h -17 l 17,-5 z m -17,0 17,-5 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8704" />
        </g>
        <g
           id="g8706">
          <path
             d="m 850,1401 h -16 l 16,-5 z m -16,0 16,-5 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8708" />
        </g>
        <g
           id="g8710">
          <path
             d="m 886,1396 h 17 v 0 z m 17,0 v 0 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8712" />
        </g>
        <g
           id="g8714">
          <path
             d="m 850,1396 h -17 l 17,-1 z m -17,0 17,-1 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8716" />
        </g>
        <g
           id="g8718">
          <path
             d="m 903,1396 h -17 l 17,-3 z m -17,0 17,-3 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8720" />
        </g>
        <g
           id="g8722">
          <path
             d="m 850,1395 h -17 l 17,-3 z m -17,0 17,-3 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8724" />
        </g>
        <g
           id="g8726">
          <path
             d="m 903,1393 h -17 l 17,-1 z m -17,0 17,-1 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8728" />
        </g>
        <g
           id="g8730">
          <path
             d="m 850,1392 h -17 l 17,-1 z m -17,0 17,-1 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8732" />
        </g>
        <g
           id="g8734">
          <path
             d="m 903,1392 h -17 l 18,-3 z m -17,0 18,-3 h -19 z m 18,-3 h -19 z m -19,0 h 19 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8736" />
        </g>
        <g
           id="g8738">
          <path
             d="m 850,1391 h -17 l 19,-3 z m -17,0 19,-3 h -21 z m 19,-3 h -21 z m -21,0 h 21 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8740" />
        </g>
        <g
           id="g8742">
          <path
             d="m 904,1389 h -19 l 20,-1 z m -19,0 20,-1 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8744" />
        </g>
        <g
           id="g8746">
          <path
             d="m 852,1388 h -21 l 23,-1 z m -21,0 23,-1 h -24 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8748" />
        </g>
        <g
           id="g8750">
          <path
             d="m 905,1388 h -22 l 25,-2 z m -22,0 25,-2 h -27 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8752" />
        </g>
        <g
           id="g8754">
          <path
             d="m 854,1387 h -24 l 26,-1 z m -24,0 26,-1 h -29 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8756" />
        </g>
        <g
           id="g8758">
          <path
             d="m 856,1386 h -29 l 29,-1 z m -29,0 29,-1 h -30 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8760" />
        </g>
        <g
           id="g8762">
          <path
             d="m 908,1386 h -27 l 28,-1 z m -27,0 28,-1 h -29 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8764" />
        </g>
        <g
           id="g8766">
          <path
             d="m 909,1385 h -29 31 z m -29,0 h 31 -33 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8768" />
        </g>
        <g
           id="g8770">
          <path
             d="m 856,1385 h -30 34 z m -30,0 h 34 -39 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8772" />
        </g>
        <g
           id="g8774">
          <path
             d="m 911,1385 h -33 34 z m -33,0 h 34 -35 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8776" />
        </g>
        <g
           id="g8778">
          <path
             d="m 912,1385 h -35 39 z m -35,0 h 39 -42 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8780" />
        </g>
        <g
           id="g8782">
          <path
             d="m 860,1385 h -39 43 z m -39,0 h 43 -44 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8784" />
        </g>
        <g
           id="g8786">
          <path
             d="m 916,1385 h -44 l 44,-4 z m -44,0 44,-4 h -44 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8788" />
        </g>
        <g
           id="g8790">
          <path
             d="m 864,1385 h -44 l 44,-4 z m -44,0 44,-4 h -44 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8792" />
        </g>
        <g
           id="g8794">
          <path
             d="m 966,1473 7,-1 h -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8796" />
        </g>
        <g
           id="g8798">
          <path
             d="m 973,1472 h -14 15 z m -14,0 h 15 -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8800" />
        </g>
        <g
           id="g8802">
          <path
             d="m 974,1472 h -17 l 22,-2 z m -17,0 22,-2 h -27 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8804" />
        </g>
        <g
           id="g8806">
          <path
             d="m 979,1470 h -27 29 z m -27,0 h 29 -31 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8808" />
        </g>
        <g
           id="g8810">
          <path
             d="m 981,1470 h -31 l 35,-3 z m -31,0 35,-3 h -40 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8812" />
        </g>
        <g
           id="g8814">
          <path
             d="m 985,1467 h -40 l 42,-1 z m -40,0 42,-1 h -44 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8816" />
        </g>
        <g
           id="g8818">
          <path
             d="m 987,1466 h -29 z m -29,0 h 29 -25 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8820" />
        </g>
        <g
           id="g8822">
          <path
             d="m 943,1466 h 15 v 0 z m 15,0 v 0 h -15 z m 0,0 h -15 z m -15,0 h 15 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8824" />
        </g>
        <g
           id="g8826">
          <path
             d="m 987,1466 h -25 l 26,-1 z m -25,0 26,-1 h -23 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8828" />
        </g>
        <g
           id="g8830">
          <path
             d="m 958,1466 h -15 l 11,-1 z m -15,0 11,-1 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8832" />
        </g>
        <g
           id="g8834">
          <path
             d="m 988,1465 h -23 l 25,-2 z m -23,0 25,-2 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8836" />
        </g>
        <g
           id="g8838">
          <path
             d="m 954,1465 h -13 l 8,-3 z m -13,0 8,-3 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8840" />
        </g>
        <g
           id="g8842">
          <path
             d="m 990,1463 h -20 l 21,-1 z m -20,0 21,-1 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8844" />
        </g>
        <g
           id="g8846">
          <path
             d="m 949,1462 h -10 l 7,-2 z m -10,0 7,-2 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8848" />
        </g>
        <g
           id="g8850">
          <path
             d="m 946,1460 h -10 l 9,-1 z m -10,0 9,-1 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8852" />
        </g>
        <g
           id="g8854">
          <path
             d="m 991,1462 h -19 l 23,-4 z m -19,0 23,-4 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8856" />
        </g>
        <g
           id="g8858">
          <path
             d="m 995,1458 h -19 l 19,-1 z m -19,0 19,-1 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8860" />
        </g>
        <g
           id="g8862">
          <path
             d="m 945,1459 h -10 l 7,-5 z m -10,0 7,-5 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8864" />
        </g>
        <g
           id="g8866">
          <path
             d="m 942,1454 h -10 l 9,-1 z m -10,0 9,-1 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8868" />
        </g>
        <g
           id="g8870">
          <path
             d="m 995,1457 h -19 l 22,-6 z m -19,0 22,-6 h -19 z m 22,-6 h -19 z m -19,0 h 19 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8872" />
        </g>
        <g
           id="g8874">
          <path
             d="m 941,1453 h -10 l 9,-4 z m -10,0 9,-4 h -11 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8876" />
        </g>
        <g
           id="g8878">
          <path
             d="m 998,1451 h -19 l 20,-4 z m -19,0 20,-4 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8880" />
        </g>
        <g
           id="g8882">
          <path
             d="m 940,1449 h -11 l 10,-4 z m -11,0 10,-4 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8884" />
        </g>
        <g
           id="g8886">
          <path
             d="m 999,1447 h -20 l 20,-3 z m -20,0 20,-3 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8888" />
        </g>
        <g
           id="g8890">
          <path
             d="m 999,1444 h -19 l 20,-2 z m -19,0 20,-2 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8892" />
        </g>
        <g
           id="g8894">
          <path
             d="m 939,1445 h -12 l 11,-3 z m -12,0 11,-3 h -11 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8896" />
        </g>
        <g
           id="g8898">
          <path
             d="m 1000,1442 h -73 l 73,-5 z m -73,0 73,-5 h -74 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8900" />
        </g>
        <g
           id="g8902">
          <path
             d="m 938,1437 h -12 l 12,-2 z m -12,0 12,-2 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8904" />
        </g>
        <g
           id="g8906">
          <path
             d="m 938,1435 h -13 l 14,-8 z m -13,0 14,-8 h -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8908" />
        </g>
        <g
           id="g8910">
          <path
             d="m 939,1427 h -14 l 15,-3 z m -14,0 15,-3 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8912" />
        </g>
        <g
           id="g8914">
          <path
             d="m 940,1424 h -15 l 16,-5 z m -15,0 16,-5 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8916" />
        </g>
        <g
           id="g8918">
          <path
             d="m 997,1416 2,-2 h -3 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8920" />
        </g>
        <g
           id="g8922">
          <path
             d="m 941,1419 h -16 l 18,-5 z m -16,0 18,-5 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8924" />
        </g>
        <g
           id="g8926">
          <path
             d="m 1000,1414 v 0 h -4 z m 0,0 h -4 3 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8928" />
        </g>
        <g
           id="g8930">
          <path
             d="m 943,1414 h -18 l 19,-2 z m -18,0 19,-2 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8932" />
        </g>
        <g
           id="g8934">
          <path
             d="m 1000,1414 h -4 l 3,-7 z m -4,0 3,-7 h -6 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8936" />
        </g>
        <g
           id="g8938">
          <path
             d="m 999,1407 h -6 l 5,-1 z m -6,0 5,-1 h -6 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8940" />
        </g>
        <g
           id="g8942">
          <path
             d="m 944,1412 h -18 l 22,-7 z m -18,0 22,-7 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8944" />
        </g>
        <g
           id="g8946">
          <path
             d="m 998,1406 h -6 l 4,-5 z m -6,0 4,-5 h -8 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8948" />
        </g>
        <g
           id="g8950">
          <path
             d="m 948,1405 h -21 l 26,-4 z m -21,0 26,-4 h -23 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8952" />
        </g>
        <g
           id="g8954">
          <path
             d="m 996,1401 h -8 l 7,-2 z m -8,0 7,-2 h -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8956" />
        </g>
        <g
           id="g8958">
          <path
             d="m 953,1401 h -23 l 28,-3 z m -23,0 28,-3 h -27 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8960" />
        </g>
        <g
           id="g8962">
          <path
             d="m 958,1398 h -27 l 28,-1 z m -27,0 28,-1 h -28 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8964" />
        </g>
        <g
           id="g8966">
          <path
             d="m 995,1399 h -9 l 7,-4 z m -9,0 7,-4 h -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8968" />
        </g>
        <g
           id="g8970">
          <path
             d="m 959,1397 h -28 l 34,-2 z m -28,0 34,-2 h -32 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8972" />
        </g>
        <g
           id="g8974">
          <path
             d="m 993,1395 h -14 z m -14,0 h 14 -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8976" />
        </g>
        <g
           id="g8978">
          <path
             d="m 933,1395 h 32 v 0 z m 32,0 v 0 h -32 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8980" />
        </g>
        <g
           id="g8982">
          <path
             d="m 993,1395 h -17 l 16,-1 z m -17,0 16,-1 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8984" />
        </g>
        <g
           id="g8986">
          <path
             d="m 965,1395 h -32 l 38,-1 z m -32,0 38,-1 h -38 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8988" />
        </g>
        <g
           id="g8990">
          <path
             d="m 992,1394 h -59 l 56,-3 z m -59,0 56,-3 h -53 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8992" />
        </g>
        <g
           id="g8994">
          <path
             d="m 989,1391 h -53 l 52,-2 z m -53,0 52,-2 h -50 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path8996" />
        </g>
        <g
           id="g8998">
          <path
             d="m 988,1389 h -50 l 46,-4 z m -50,0 46,-4 h -42 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9000" />
        </g>
        <g
           id="g9002">
          <path
             d="m 984,1385 h -42 l 41,-1 z m -42,0 41,-1 h -40 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9004" />
        </g>
        <g
           id="g9006">
          <path
             d="m 983,1384 h -40 l 35,-3 z m -40,0 35,-3 h -29 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9008" />
        </g>
        <g
           id="g9010">
          <path
             d="m 978,1381 h -29 28 z m -29,0 h 28 -27 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9012" />
        </g>
        <g
           id="g9014">
          <path
             d="m 977,1381 h -27 l 21,-2 z m -27,0 21,-2 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9016" />
        </g>
        <g
           id="g9018">
          <path
             d="m 956,1379 h 1 14 z m 1,0 h 14 l -7,-1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9020" />
        </g>
        <g
           id="g9022">
          <path
             d="m 956,1379 h 15 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9024" />
        </g>
        <g
           id="g9026">
          <path
             d="m 1131,1516 h 2 -8 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9028" />
        </g>
        <g
           id="g9030">
          <path
             d="m 1133,1516 h -8 11 z m -8,0 h 11 -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9032" />
        </g>
        <g
           id="g9034">
          <path
             d="m 1136,1516 h -12 l 21,-2 z m -12,0 21,-2 h -32 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9036" />
        </g>
        <g
           id="g9038">
          <path
             d="m 1146,1514 v 0 h -33 z m 0,0 h -33 32 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9040" />
        </g>
        <g
           id="g9042">
          <path
             d="m 1176,1516 h -4 l 4,-5 z m -4,0 4,-5 h -6 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9044" />
        </g>
        <g
           id="g9046">
          <path
             d="m 1146,1514 h -33 l 43,-4 z m -33,0 43,-4 h -53 z m 43,-4 h -53 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9048" />
        </g>
        <g
           id="g9050">
          <path
             d="m 1103,1510 h 53 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9052" />
        </g>
        <g
           id="g9054">
          <path
             d="m 1156,1510 h -54 l 56,-1 z m -54,0 56,-1 h -58 z m 56,-1 h -58 z m -58,0 h 58 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9056" />
        </g>
        <g
           id="g9058">
          <path
             d="m 1127,1509 v 0 h -27 z m 0,0 h -27 36 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9060" />
        </g>
        <g
           id="g9062">
          <path
             d="m 1158,1509 h -22 23 z m -22,0 h 23 -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9064" />
        </g>
        <g
           id="g9066">
          <path
             d="m 1159,1509 h -22 l 23,-1 z m -22,0 23,-1 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9068" />
        </g>
        <g
           id="g9070">
          <path
             d="m 1176,1511 h -6 l 6,-3 z m -6,0 6,-3 h -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9072" />
        </g>
        <g
           id="g9074">
          <path
             d="m 1127,1509 h -27 l 19,-1 z m -27,0 19,-1 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9076" />
        </g>
        <g
           id="g9078">
          <path
             d="m 1160,1508 h -19 21 z m -19,0 h 21 -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9080" />
        </g>
        <g
           id="g9082">
          <path
             d="m 1176,1508 h -9 l 9,-1 z m -9,0 9,-1 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9084" />
        </g>
        <g
           id="g9086">
          <path
             d="m 1162,1508 h -18 l 20,-1 z m -18,0 20,-1 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9088" />
        </g>
        <g
           id="g9090">
          <path
             d="m 1119,1508 h -21 l 14,-3 z m -21,0 14,-3 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9092" />
        </g>
        <g
           id="g9094">
          <path
             d="m 1176,1507 h -30 l 30,-3 z m -30,0 30,-3 h -23 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9096" />
        </g>
        <g
           id="g9098">
          <path
             d="m 1112,1505 h -19 l 18,-1 z m -19,0 18,-1 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9100" />
        </g>
        <g
           id="g9102">
          <path
             d="m 1111,1504 h -20 l 14,-3 z m -20,0 14,-3 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9104" />
        </g>
        <g
           id="g9106">
          <path
             d="m 1176,1504 h -23 l 24,-5 z m -23,0 24,-5 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9108" />
        </g>
        <g
           id="g9110">
          <path
             d="m 1105,1501 h -17 l 12,-5 z m -17,0 12,-5 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9112" />
        </g>
        <g
           id="g9114">
          <path
             d="m 1100,1496 h -18 l 18,-1 z m -18,0 18,-1 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9116" />
        </g>
        <g
           id="g9118">
          <path
             d="m 1177,1499 h -17 l 17,-7 z m -17,0 17,-7 h -11 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9120" />
        </g>
        <g
           id="g9122">
          <path
             d="m 1100,1495 h -18 l 13,-7 z m -18,0 13,-7 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9124" />
        </g>
        <g
           id="g9126">
          <path
             d="m 1095,1488 h -19 l 18,-2 z m -19,0 18,-2 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9128" />
        </g>
        <g
           id="g9130">
          <path
             d="m 1177,1492 h -11 l 12,-9 z m -11,0 12,-9 h -7 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9132" />
        </g>
        <g
           id="g9134">
          <path
             d="m 1094,1486 h -19 l 16,-7 z m -19,0 16,-7 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9136" />
        </g>
        <g
           id="g9138">
          <path
             d="m 1091,1479 h -20 l 18,-4 z m -20,0 18,-4 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9140" />
        </g>
        <g
           id="g9142">
          <path
             d="m 1178,1483 h -7 l 8,-12 z m -7,0 8,-12 h -3 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9144" />
        </g>
        <g
           id="g9146">
          <path
             d="m 1089,1475 h -20 l 19,-6 z m -20,0 19,-6 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9148" />
        </g>
        <g
           id="g9150">
          <path
             d="m 1088,1469 h -21 l 20,-6 z m -21,0 20,-6 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9152" />
        </g>
        <g
           id="g9154">
          <path
             d="m 1087,1463 h -22 l 21,-5 z m -22,0 21,-5 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9156" />
        </g>
        <g
           id="g9158">
          <path
             d="m 1086,1458 h -22 l 21,-8 z m -22,0 21,-8 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9160" />
        </g>
        <g
           id="g9162">
          <path
             d="m 1085,1450 h -22 l 22,-5 z m -22,0 22,-5 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9164" />
        </g>
        <g
           id="g9166">
          <path
             d="m 1085,1445 h -22 l 22,-2 z m -22,0 22,-2 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9168" />
        </g>
        <g
           id="g9170">
          <path
             d="m 1085,1443 h -22 l 23,-8 z m -22,0 23,-8 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9172" />
        </g>
        <g
           id="g9174">
          <path
             d="m 1086,1435 h -22 l 22,-1 z m -22,0 22,-1 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9176" />
        </g>
        <g
           id="g9178">
          <path
             d="m 1086,1434 h -22 l 23,-10 z m -22,0 23,-10 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9180" />
        </g>
        <g
           id="g9182">
          <path
             d="m 1087,1424 h -21 l 23,-5 z m -21,0 23,-5 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9184" />
        </g>
        <g
           id="g9186">
          <path
             d="m 1089,1419 h -22 l 23,-4 z m -22,0 23,-4 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9188" />
        </g>
        <g
           id="g9190">
          <path
             d="m 1179,1414 3,-2 h -5 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9192" />
        </g>
        <g
           id="g9194">
          <path
             d="m 1090,1415 h -21 l 25,-7 z m -21,0 25,-7 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9196" />
        </g>
        <g
           id="g9198">
          <path
             d="m 1094,1408 h -21 l 22,-2 z m -21,0 22,-2 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9200" />
        </g>
        <g
           id="g9202">
          <path
             d="m 1182,1412 h -5 v -7 z m -5,0 v -7 h -5 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9204" />
        </g>
        <g
           id="g9206">
          <path
             d="m 1095,1406 h -21 l 24,-3 z m -21,0 24,-3 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9208" />
        </g>
        <g
           id="g9210">
          <path
             d="m 1177,1405 h -5 l 3,-4 z m -5,0 3,-4 h -7 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9212" />
        </g>
        <g
           id="g9214">
          <path
             d="m 1098,1403 h -22 l 23,-2 z m -22,0 23,-2 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9216" />
        </g>
        <g
           id="g9218">
          <path
             d="m 1099,1401 h -21 l 24,-2 z m -21,0 24,-2 h -23 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9220" />
        </g>
        <g
           id="g9222">
          <path
             d="m 1175,1401 h -7 l 4,-3 z m -7,0 4,-3 h -7 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9224" />
        </g>
        <g
           id="g9226">
          <path
             d="m 1102,1399 h -23 l 26,-4 z m -23,0 26,-4 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9228" />
        </g>
        <g
           id="g9230">
          <path
             d="m 1172,1398 h -7 l 2,-5 z m -7,0 2,-5 h -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9232" />
        </g>
        <g
           id="g9234">
          <path
             d="m 1167,1393 h -9 l 9,-1 z m -9,0 9,-1 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9236" />
        </g>
        <g
           id="g9238">
          <path
             d="m 1105,1395 h -22 l 29,-3 z m -22,0 29,-3 h -26 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9240" />
        </g>
        <g
           id="g9242">
          <path
             d="m 1112,1392 h -26 l 27,-1 z m -26,0 27,-1 h -26 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9244" />
        </g>
        <g
           id="g9246">
          <path
             d="m 1167,1392 h -10 l 6,-2 z m -10,0 6,-2 h -11 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9248" />
        </g>
        <g
           id="g9250">
          <path
             d="m 1113,1391 h -26 l 34,-3 z m -26,0 34,-3 h -30 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9252" />
        </g>
        <g
           id="g9254">
          <path
             d="m 1163,1390 h -11 l 8,-2 z m -11,0 8,-2 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9256" />
        </g>
        <g
           id="g9258">
          <path
             d="m 1160,1388 h -15 l 14,-1 z m -15,0 14,-1 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9260" />
        </g>
        <g
           id="g9262">
          <path
             d="m 1121,1388 h -30 l 38,-1 z m -30,0 38,-1 h -36 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9264" />
        </g>
        <g
           id="g9266">
          <path
             d="m 1159,1387 h -20 z m -20,0 h 20 -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9268" />
        </g>
        <g
           id="g9270">
          <path
             d="m 1138,1387 v 0 h -45 z m 0,0 h -45 36 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9272" />
        </g>
        <g
           id="g9274">
          <path
             d="m 1159,1387 h -66 l 65,-1 z m -66,0 65,-1 h -64 z m 65,-1 h -64 1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9276" />
        </g>
        <g
           id="g9278">
          <path
             d="m 1094,1386 h 64 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9280" />
        </g>
        <g
           id="g9282">
          <path
             d="m 1158,1386 h -63 l 55,-4 z m -63,0 55,-4 h -47 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9284" />
        </g>
        <g
           id="g9286">
          <path
             d="m 1150,1382 h -47 l 45,-1 z m -47,0 45,-1 h -42 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9288" />
        </g>
        <g
           id="g9290">
          <path
             d="m 1148,1381 h -42 l 34,-2 z m -42,0 34,-2 h -27 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9292" />
        </g>
        <g
           id="g9294">
          <path
             d="m 1140,1379 h -27 24 z m -27,0 h 24 -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9296" />
        </g>
        <g
           id="g9298">
          <path
             d="m 1137,1379 h -19 l 13,-1 z m -19,0 13,-1 h -8 z m 13,-1 h -8 5 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9300" />
        </g>
        <g
           id="g9302">
          <path
             d="m 1123,1378 h 8 v 0 z m 8,0 v 0 h -8 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9304" />
        </g>
        <g
           id="g9306">
          <path
             d="m 1226,1473 h -5 l 5,-11 z m -5,0 5,-11 h -32 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9308" />
        </g>
        <g
           id="g9310">
          <path
             d="m 1226,1462 h -32 l 32,-2 z m -32,0 32,-2 h -31 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9312" />
        </g>
        <g
           id="g9314">
          <path
             d="m 1196,1459 h 1 l -1,-1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9316" />
        </g>
        <g
           id="g9318">
          <path
             d="m 1226,1460 h -24 l 24,-1 z m -24,0 24,-1 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9320" />
        </g>
        <g
           id="g9322">
          <path
             d="m 1202,1460 h -7 l 2,-1 z m -7,0 2,-1 h -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9324" />
        </g>
        <g
           id="g9326">
          <path
             d="m 1226,1459 h -20 l 20,-2 z m -20,0 20,-2 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9328" />
        </g>
        <g
           id="g9330">
          <path
             d="m 1226,1457 h -18 l 18,-3 z m -18,0 18,-3 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9332" />
        </g>
        <g
           id="g9334">
          <path
             d="m 1226,1454 h -17 l 17,-2 z m -17,0 17,-2 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9336" />
        </g>
        <g
           id="g9338">
          <path
             d="m 1226,1452 h -17 l 17,-5 z m -17,0 17,-5 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9340" />
        </g>
        <g
           id="g9342">
          <path
             d="m 1226,1447 h -17 l 17,-5 z m -17,0 17,-5 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9344" />
        </g>
        <g
           id="g9346">
          <path
             d="m 1226,1442 h -17 l 17,-6 z m -17,0 17,-6 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9348" />
        </g>
        <g
           id="g9350">
          <path
             d="m 1226,1436 h -17 l 17,-35 z m -17,0 17,-35 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9352" />
        </g>
        <g
           id="g9354">
          <path
             d="m 1226,1401 h -17 l 17,-5 z m -17,0 17,-5 h -17 z m 17,-5 h -17 z m -17,0 h 17 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9356" />
        </g>
        <g
           id="g9358">
          <path
             d="m 1226,1396 h -17 l 17,-4 z m -17,0 17,-4 h -17 z m 17,-4 h -17 z m -17,0 h 17 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9360" />
        </g>
        <g
           id="g9362">
          <path
             d="m 1226,1392 h -17 l 19,-4 z m -17,0 19,-4 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9364" />
        </g>
        <g
           id="g9366">
          <path
             d="m 1229,1388 v 0 h -22 z m 0,0 h -22 21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9368" />
        </g>
        <g
           id="g9370">
          <path
             d="m 1229,1388 h -22 l 25,-3 z m -22,0 25,-3 h -29 z m 25,-3 h -29 z m -29,0 h 29 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9372" />
        </g>
        <g
           id="g9374">
          <path
             d="m 1232,1385 h -29 32 z m -29,0 h 32 -35 z m 32,0 h -35 z m -35,0 h 35 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9376" />
        </g>
        <g
           id="g9378">
          <path
             d="m 1235,1385 h -35 39 z m -35,0 h 39 -43 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9380" />
        </g>
        <g
           id="g9382">
          <path
             d="m 1239,1385 h -43 l 43,-4 z m -43,0 43,-4 h -43 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9384" />
        </g>
        <g
           id="g9386">
          <path
             d="m 1276,1500 h -3 l 3,-7 z m -3,0 3,-7 h -5 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9388" />
        </g>
        <g
           id="g9390">
          <path
             d="m 1276,1493 h -5 l 5,-5 z m -5,0 5,-5 h -8 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9392" />
        </g>
        <g
           id="g9394">
          <path
             d="m 1276,1488 h -8 l 8,-4 z m -8,0 8,-4 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9396" />
        </g>
        <g
           id="g9398">
          <path
             d="m 1276,1484 h -10 l 10,-4 z m -10,0 10,-4 h -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9400" />
        </g>
        <g
           id="g9402">
          <path
             d="m 1276,1480 h -14 l 14,-8 z m -14,0 14,-8 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9404" />
        </g>
        <g
           id="g9406">
          <path
             d="m 1276,1472 h -22 l 22,-2 z m -22,0 22,-2 h -24 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9408" />
        </g>
        <g
           id="g9410">
          <path
             d="m 1297,1470 h -45 l 45,-3 z m -45,0 45,-3 h -51 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9412" />
        </g>
        <g
           id="g9414">
          <path
             d="m 1297,1467 h -51 l 51,-4 z m -51,0 51,-4 h -51 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9416" />
        </g>
        <g
           id="g9418">
          <path
             d="m 1276,1463 h -16 l 16,-57 z m -16,0 16,-57 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9420" />
        </g>
        <g
           id="g9422">
          <path
             d="m 1276,1406 h -16 l 17,-3 z m -16,0 17,-3 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9424" />
        </g>
        <g
           id="g9426">
          <path
             d="m 1277,1403 h -17 l 17,-5 z m -17,0 17,-5 h -17 z m 17,-5 h -17 z m -17,0 h 17 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9428" />
        </g>
        <g
           id="g9430">
          <path
             d="m 1300,1399 h -4 l 3,-4 z m -4,0 3,-4 h -5 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9432" />
        </g>
        <g
           id="g9434">
          <path
             d="m 1277,1398 h -17 l 19,-4 z m -17,0 19,-4 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9436" />
        </g>
        <g
           id="g9438">
          <path
             d="m 1279,1394 h -18 l 19,-1 z m -18,0 19,-1 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9440" />
        </g>
        <g
           id="g9442">
          <path
             d="m 1299,1395 h -5 l 4,-2 z m -5,0 4,-2 h -6 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9444" />
        </g>
        <g
           id="g9446">
          <path
             d="m 1297,1393 v 0 h -5 z m 0,0 h -5 6 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9448" />
        </g>
        <g
           id="g9450">
          <path
             d="m 1280,1393 h -19 l 21,-1 z m -19,0 21,-1 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9452" />
        </g>
        <g
           id="g9454">
          <path
             d="m 1297,1393 h -5 l 4,-2 z m -5,0 4,-2 h -8 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9456" />
        </g>
        <g
           id="g9458">
          <path
             d="m 1282,1392 h -20 l 21,-1 z m -20,0 21,-1 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9460" />
        </g>
        <g
           id="g9462">
          <path
             d="m 1296,1391 h -8 z m -8,0 h 8 -11 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9464" />
        </g>
        <g
           id="g9466">
          <path
             d="m 1285,1391 v 0 h -23 z m 0,0 h -23 21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9468" />
        </g>
        <g
           id="g9470">
          <path
             d="m 1296,1391 h -34 l 33,-2 z m -34,0 33,-2 h -32 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9472" />
        </g>
        <g
           id="g9474">
          <path
             d="m 1295,1389 h -32 l 30,-2 z m -32,0 30,-2 h -30 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9476" />
        </g>
        <g
           id="g9478">
          <path
             d="m 1293,1387 h -30 l 28,-2 z m -30,0 28,-2 h -26 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9480" />
        </g>
        <g
           id="g9482">
          <path
             d="m 1291,1385 h -26 l 23,-2 z m -26,0 23,-2 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9484" />
        </g>
        <g
           id="g9486">
          <path
             d="m 1288,1383 h -20 l 19,-1 z m -20,0 19,-1 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9488" />
        </g>
        <g
           id="g9490">
          <path
             d="m 1268,1382 5,-2 h 8 z m 5,-2 h 8 -2 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9492" />
        </g>
        <g
           id="g9494">
          <path
             d="m 1268,1382 h 19 l -6,-2 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9496" />
        </g>
        <g
           id="g9498">
          <path
             d="m 1398,1470 h -29 l 29,-3 z m -29,0 29,-3 h -29 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9500" />
        </g>
        <g
           id="g9502">
          <path
             d="m 1342,1470 h -41 l 41,-3 z m -41,0 41,-3 h -41 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9504" />
        </g>
        <g
           id="g9506">
          <path
             d="m 1398,1467 h -29 28 z m -29,0 h 28 -24 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9508" />
        </g>
        <g
           id="g9510">
          <path
             d="m 1397,1467 h -24 l 22,-1 z m -24,0 22,-1 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9512" />
        </g>
        <g
           id="g9514">
          <path
             d="m 1395,1466 h -20 19 z m -20,0 h 19 -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9516" />
        </g>
        <g
           id="g9518">
          <path
             d="m 1340,1467 h -39 l 34,-1 z m -39,0 34,-1 h -31 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9520" />
        </g>
        <g
           id="g9522">
          <path
             d="m 1335,1466 h -31 l 30,-1 z m -31,0 30,-1 h -27 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9524" />
        </g>
        <g
           id="g9526">
          <path
             d="m 1394,1466 h -18 l 16,-2 z m -18,0 16,-2 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9528" />
        </g>
        <g
           id="g9530">
          <path
             d="m 1392,1464 h -15 l 14,-1 z m -15,0 14,-1 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9532" />
        </g>
        <g
           id="g9534">
          <path
             d="m 1334,1465 h -27 l 25,-2 z m -27,0 25,-2 h -23 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9536" />
        </g>
        <g
           id="g9538">
          <path
             d="m 1332,1463 h -23 l 23,-1 z m -23,0 23,-1 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9540" />
        </g>
        <g
           id="g9542">
          <path
             d="m 1391,1463 h -13 l 11,-1 z m -13,0 11,-1 h -11 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9544" />
        </g>
        <g
           id="g9546">
          <path
             d="m 1332,1462 h -22 l 22,-1 z m -22,0 22,-1 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9548" />
        </g>
        <g
           id="g9550">
          <path
             d="m 1332,1461 h -21 l 21,-1 z m -21,0 21,-1 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9552" />
        </g>
        <g
           id="g9554">
          <path
             d="m 1389,1462 h -11 l 10,-2 z m -11,0 10,-2 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9556" />
        </g>
        <g
           id="g9558">
          <path
             d="m 1332,1460 h -21 l 21,-2 z m -21,0 21,-2 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9560" />
        </g>
        <g
           id="g9562">
          <path
             d="m 1332,1458 h -19 l 19,-1 z m -19,0 19,-1 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9564" />
        </g>
        <g
           id="g9566">
          <path
             d="m 1388,1460 h -10 l 9,-3 z m -10,0 9,-3 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9568" />
        </g>
        <g
           id="g9570">
          <path
             d="m 1332,1457 h -19 l 20,-3 z m -19,0 20,-3 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9572" />
        </g>
        <g
           id="g9574">
          <path
             d="m 1387,1457 h -10 l 8,-3 z m -10,0 8,-3 h -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9576" />
        </g>
        <g
           id="g9578">
          <path
             d="m 1385,1454 h -9 l 9,-1 z m -9,0 9,-1 h -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9580" />
        </g>
        <g
           id="g9582">
          <path
             d="m 1333,1454 h -18 l 19,-2 z m -18,0 19,-2 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9584" />
        </g>
        <g
           id="g9586">
          <path
             d="m 1385,1453 h -9 l 7,-3 z m -9,0 7,-3 h -8 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9588" />
        </g>
        <g
           id="g9590">
          <path
             d="m 1334,1452 h -17 l 18,-2 z m -17,0 18,-2 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9592" />
        </g>
        <g
           id="g9594">
          <path
             d="m 1383,1450 h -8 l -10,-46 z m -8,0 -10,-46 h -8 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9596" />
        </g>
        <g
           id="g9598">
          <path
             d="m 1335,1450 h -17 l 39,-46 z m -17,0 39,-46 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9600" />
        </g>
        <g
           id="g9602">
          <path
             d="m 1365,1404 h -26 l 18,-19 z m -26,0 18,-19 h -8 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9604" />
        </g>
        <g
           id="g9606">
          <path
             d="m 1357,1385 h -8 l 2,-16 z m -8,0 2,-16 h -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9608" />
        </g>
        <g
           id="g9610">
          <path
             d="m 1351,1369 h -9 l 7,-5 z m -9,0 7,-5 h -9 z m 7,-5 h -9 z m -9,0 h 9 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9612" />
        </g>
        <g
           id="g9614">
          <path
             d="m 1349,1364 h -9 l 7,-3 z m -9,0 7,-3 h -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9616" />
        </g>
        <g
           id="g9618">
          <path
             d="m 1317,1358 h 1 -6 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9620" />
        </g>
        <g
           id="g9622">
          <path
             d="m 1347,1361 h -9 l 7,-4 z m -9,0 7,-4 h -11 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9624" />
        </g>
        <g
           id="g9626">
          <path
             d="m 1318,1358 h -6 l 11,-2 z m -6,0 11,-2 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9628" />
        </g>
        <g
           id="g9630">
          <path
             d="m 1345,1357 h -11 l 11,-1 z m -11,0 11,-1 h -11 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9632" />
        </g>
        <g
           id="g9634">
          <path
             d="m 1323,1356 h -13 15 z m -13,0 h 15 -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9636" />
        </g>
        <g
           id="g9638">
          <path
             d="m 1325,1356 h -17 l 17,-1 z m -17,0 17,-1 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9640" />
        </g>
        <g
           id="g9642">
          <path
             d="m 1327,1355 v 0 h -19 z m 0,0 h -19 17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9644" />
        </g>
        <g
           id="g9646">
          <path
             d="m 1345,1356 h -11 l 10,-1 z m -11,0 10,-1 h -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9648" />
        </g>
        <g
           id="g9650">
          <path
             d="m 1327,1355 h -19 22 z m -19,0 h 22 -23 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9652" />
        </g>
        <g
           id="g9654">
          <path
             d="m 1344,1355 h -37 l 35,-3 z m -37,0 35,-3 h -36 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9656" />
        </g>
        <g
           id="g9658">
          <path
             d="m 1342,1352 h -36 l 35,-1 z m -36,0 35,-1 h -35 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9660" />
        </g>
        <g
           id="g9662">
          <path
             d="m 1341,1351 h -35 l 31,-4 z m -35,0 31,-4 h -31 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9664" />
        </g>
        <g
           id="g9666">
          <path
             d="m 1337,1347 h -31 l 30,-1 z m -31,0 30,-1 h -30 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9668" />
        </g>
        <g
           id="g9670">
          <path
             d="m 1336,1346 h -30 l 25,-4 z m -30,0 25,-4 h -23 z m 25,-4 h -23 1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9672" />
        </g>
        <g
           id="g9674">
          <path
             d="m 1308,1342 h 23 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9676" />
        </g>
        <g
           id="g9678">
          <path
             d="m 1331,1342 h -22 l 16,-3 z m -22,0 16,-3 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9680" />
        </g>
        <g
           id="g9682">
          <path
             d="m 1324,1339 v 0 h -11 z m 0,0 h -11 12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9684" />
        </g>
        <g
           id="g9686">
          <path
             d="m 1313,1339 3,-1 h 5 z m 3,-1 h 5 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9688" />
        </g>
        <g
           id="g9690">
          <path
             d="m 1313,1339 h 11 l -3,-1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9692" />
        </g>
        <g
           id="g9694">
          <path
             d="m 1499,1473 5,-1 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9696" />
        </g>
        <g
           id="g9698">
          <path
             d="m 1504,1472 h -12 l 19,-1 z m -12,0 19,-1 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9700" />
        </g>
        <g
           id="g9702">
          <path
             d="m 1511,1471 h -22 24 z m -22,0 h 24 -27 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9704" />
        </g>
        <g
           id="g9706">
          <path
             d="m 1513,1471 h -27 l 33,-3 z m -27,0 33,-3 h -40 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9708" />
        </g>
        <g
           id="g9710">
          <path
             d="m 1519,1468 h -40 l 42,-1 z m -40,0 42,-1 h -43 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9712" />
        </g>
        <g
           id="g9714">
          <path
             d="m 1521,1467 h -43 l 44,-1 z m -43,0 44,-1 h -45 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9716" />
        </g>
        <g
           id="g9718">
          <path
             d="m 1522,1466 h -26 27 z m -26,0 h 27 -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9720" />
        </g>
        <g
           id="g9722">
          <path
             d="m 1496,1466 h -19 13 z m -19,0 h 13 -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9724" />
        </g>
        <g
           id="g9726">
          <path
             d="m 1490,1466 h -14 l 11,-2 z m -14,0 11,-2 h -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9728" />
        </g>
        <g
           id="g9730">
          <path
             d="m 1523,1466 h -21 l 23,-2 z m -21,0 23,-2 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9732" />
        </g>
        <g
           id="g9734">
          <path
             d="m 1487,1464 h -14 l 11,-1 z m -14,0 11,-1 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9736" />
        </g>
        <g
           id="g9738">
          <path
             d="m 1525,1464 h -18 l 23,-4 z m -18,0 23,-4 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9740" />
        </g>
        <g
           id="g9742">
          <path
             d="m 1530,1460 h -19 l 19,-1 z m -19,0 19,-1 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9744" />
        </g>
        <g
           id="g9746">
          <path
             d="m 1484,1463 h -12 l 9,-4 z m -12,0 9,-4 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9748" />
        </g>
        <g
           id="g9750">
          <path
             d="m 1530,1459 h -18 l 19,-2 z m -18,0 19,-2 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9752" />
        </g>
        <g
           id="g9754">
          <path
             d="m 1481,1459 h -13 l 12,-2 z m -13,0 12,-2 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9756" />
        </g>
        <g
           id="g9758">
          <path
             d="m 1531,1457 h -17 l 20,-3 z m -17,0 20,-3 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9760" />
        </g>
        <g
           id="g9762">
          <path
             d="m 1480,1457 h -13 l 10,-5 z m -13,0 10,-5 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9764" />
        </g>
        <g
           id="g9766">
          <path
             d="m 1534,1454 h -18 l 20,-3 z m -18,0 20,-3 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9768" />
        </g>
        <g
           id="g9770">
          <path
             d="m 1477,1452 h -13 l 12,-3 z m -13,0 12,-3 h -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9772" />
        </g>
        <g
           id="g9774">
          <path
             d="m 1476,1449 h -14 l 13,-4 z m -14,0 13,-4 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9776" />
        </g>
        <g
           id="g9778">
          <path
             d="m 1536,1451 h -19 l 22,-7 z m -19,0 22,-7 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9780" />
        </g>
        <g
           id="g9782">
          <path
             d="m 1539,1444 h -19 l 20,-3 z m -19,0 20,-3 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9784" />
        </g>
        <g
           id="g9786">
          <path
             d="m 1475,1445 h -15 l 14,-8 z m -15,0 14,-8 h -16 z m 14,-8 h -16 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9788" />
        </g>
        <g
           id="g9790">
          <path
             d="m 1458,1437 h 16 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9792" />
        </g>
        <g
           id="g9794">
          <path
             d="m 1474,1437 h -17 l 17,-3 z m -17,0 17,-3 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9796" />
        </g>
        <g
           id="g9798">
          <path
             d="m 1540,1441 h -19 l 21,-7 z m -19,0 21,-7 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9800" />
        </g>
        <g
           id="g9802">
          <path
             d="m 1542,1434 h -19 l 19,-3 z m -19,0 19,-3 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9804" />
        </g>
        <g
           id="g9806">
          <path
             d="m 1474,1434 h -17 l 17,-5 z m -17,0 17,-5 h -18 z m 17,-5 h -18 z m -18,0 h 18 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9808" />
        </g>
        <g
           id="g9810">
          <path
             d="m 1542,1431 h -19 l 19,-4 z m -19,0 19,-4 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9812" />
        </g>
        <g
           id="g9814">
          <path
             d="m 1474,1429 h -18 l 19,-3 z m -18,0 19,-3 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9816" />
        </g>
        <g
           id="g9818">
          <path
             d="m 1542,1427 h -18 l 18,-4 z m -18,0 18,-4 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9820" />
        </g>
        <g
           id="g9822">
          <path
             d="m 1542,1423 h -18 l 18,-2 z m -18,0 18,-2 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9824" />
        </g>
        <g
           id="g9826">
          <path
             d="m 1475,1426 h -19 l 19,-5 z m -19,0 19,-5 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9828" />
        </g>
        <g
           id="g9830">
          <path
             d="m 1475,1421 h -19 l 19,-2 z m -19,0 19,-2 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9832" />
        </g>
        <g
           id="g9834">
          <path
             d="m 1542,1421 h -18 l 17,-6 z m -18,0 17,-6 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9836" />
        </g>
        <g
           id="g9838">
          <path
             d="m 1541,1415 h -17 l 15,-4 z m -17,0 15,-4 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9840" />
        </g>
        <g
           id="g9842">
          <path
             d="m 1475,1419 h -19 l 21,-8 z m -19,0 21,-8 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9844" />
        </g>
        <g
           id="g9846">
          <path
             d="m 1477,1411 h -19 l 19,-1 z m -19,0 19,-1 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9848" />
        </g>
        <g
           id="g9850">
          <path
             d="m 1539,1411 h -15 l 14,-3 z m -15,0 14,-3 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9852" />
        </g>
        <g
           id="g9854">
          <path
             d="m 1538,1408 h -15 l 13,-5 z m -15,0 13,-5 h -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9856" />
        </g>
        <g
           id="g9858">
          <path
             d="m 1477,1410 h -19 l 23,-9 z m -19,0 23,-9 h -19 z m 23,-9 h -19 z m -19,0 h 19 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9860" />
        </g>
        <g
           id="g9862">
          <path
             d="m 1536,1403 h -14 l 13,-3 z m -14,0 13,-3 h -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9864" />
        </g>
        <g
           id="g9866">
          <path
             d="m 1535,1400 h -14 l 11,-4 z m -14,0 11,-4 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9868" />
        </g>
        <g
           id="g9870">
          <path
             d="m 1481,1401 h -19 l 23,-7 z m -19,0 23,-7 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9872" />
        </g>
        <g
           id="g9874">
          <path
             d="m 1532,1396 h -12 l 10,-3 z m -12,0 10,-3 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9876" />
        </g>
        <g
           id="g9878">
          <path
             d="m 1485,1394 h -18 l 20,-2 z m -18,0 20,-2 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9880" />
        </g>
        <g
           id="g9882">
          <path
             d="m 1530,1393 h -12 l 11,-1 z m -12,0 11,-1 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9884" />
        </g>
        <g
           id="g9886">
          <path
             d="m 1487,1392 h -19 l 23,-3 z m -19,0 23,-3 h -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9888" />
        </g>
        <g
           id="g9890">
          <path
             d="m 1529,1392 h -12 l 9,-4 z m -12,0 9,-4 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9892" />
        </g>
        <g
           id="g9894">
          <path
             d="m 1526,1388 h -13 12 z m -13,0 h 12 -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9896" />
        </g>
        <g
           id="g9898">
          <path
             d="m 1525,1388 h -13 l 11,-2 z m -13,0 11,-2 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9900" />
        </g>
        <g
           id="g9902">
          <path
             d="m 1491,1389 h -19 l 25,-3 z m -19,0 25,-3 h -22 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9904" />
        </g>
        <g
           id="g9906">
          <path
             d="m 1523,1386 h -15 l 13,-1 z m -15,0 13,-1 h -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9908" />
        </g>
        <g
           id="g9910">
          <path
             d="m 1497,1386 h -22 l 28,-1 z m -22,0 28,-1 h -28 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9912" />
        </g>
        <g
           id="g9914">
          <path
             d="m 1521,1385 h -46 45 z m -46,0 h 45 -44 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9916" />
        </g>
        <g
           id="g9918">
          <path
             d="m 1520,1385 h -44 l 43,-1 z m -44,0 43,-1 h -41 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9920" />
        </g>
        <g
           id="g9922">
          <path
             d="m 1519,1384 h -41 l 35,-3 z m -41,0 35,-3 h -29 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9924" />
        </g>
        <g
           id="g9926">
          <path
             d="m 1513,1381 h -29 l 25,-1 z m -29,0 25,-1 h -23 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9928" />
        </g>
        <g
           id="g9930">
          <path
             d="m 1486,1380 7,-1 h 13 z m 7,-1 h 13 l -8,-1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9932" />
        </g>
        <g
           id="g9934">
          <path
             d="m 1486,1380 h 23 l -3,-1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9936" />
        </g>
        <g
           id="g9938">
          <path
             d="m 1606,1526 h 4 -7 z m 4,0 h -7 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9940" />
        </g>
        <g
           id="g9942">
          <path
             d="m 1603,1526 h 7 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9944" />
        </g>
        <g
           id="g9946">
          <path
             d="m 1610,1526 h -8 l 13,-1 z m -8,0 13,-1 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9948" />
        </g>
        <g
           id="g9950">
          <path
             d="m 1615,1525 h -15 l 19,-1 z m -15,0 19,-1 h -24 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9952" />
        </g>
        <g
           id="g9954">
          <path
             d="m 1619,1524 h -24 l 24,-1 z m -24,0 24,-1 h -25 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9956" />
        </g>
        <g
           id="g9958">
          <path
             d="m 1619,1523 h -25 l 23,-5 z m -25,0 23,-5 h -32 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9960" />
        </g>
        <g
           id="g9962">
          <path
             d="m 1617,1518 h -32 l 31,-3 z m -32,0 31,-3 h -33 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9964" />
        </g>
        <g
           id="g9966">
          <path
             d="m 1616,1515 h -16 z m -16,0 h 16 -11 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9968" />
        </g>
        <g
           id="g9970">
          <path
             d="m 1583,1515 h 17 v 0 z m 17,0 v 0 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9972" />
        </g>
        <g
           id="g9974">
          <path
             d="m 1616,1515 h -11 z m -11,0 h 11 -6 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9976" />
        </g>
        <g
           id="g9978">
          <path
             d="m 1600,1515 h -17 l 12,-1 z m -17,0 12,-1 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9980" />
        </g>
        <g
           id="g9982">
          <path
             d="m 1610,1515 3,-2 h 3 z m 3,-2 h 3 l -1,-1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9984" />
        </g>
        <g
           id="g9986">
          <path
             d="m 1610,1515 h 6 v -2 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9988" />
        </g>
        <g
           id="g9990">
          <path
             d="m 1595,1514 h -13 l 9,-4 z m -13,0 9,-4 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9992" />
        </g>
        <g
           id="g9994">
          <path
             d="m 1591,1510 h -12 l 12,-1 z m -12,0 12,-1 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path9996" />
        </g>
        <g
           id="g9998">
          <path
             d="m 1591,1509 h -13 l 10,-4 z m -13,0 10,-4 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10000" />
        </g>
        <g
           id="g10002">
          <path
             d="m 1588,1505 h -12 l 10,-5 z m -12,0 10,-5 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10004" />
        </g>
        <g
           id="g10006">
          <path
             d="m 1586,1500 h -13 l 12,-2 z m -13,0 12,-2 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10008" />
        </g>
        <g
           id="g10010">
          <path
             d="m 1585,1498 h -13 l 12,-8 z m -13,0 12,-8 h -14 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10012" />
        </g>
        <g
           id="g10014">
          <path
             d="m 1584,1490 h -14 l 13,-1 z m -14,0 13,-1 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10016" />
        </g>
        <g
           id="g10018">
          <path
             d="m 1583,1489 h -13 l 12,-9 z m -13,0 12,-9 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10020" />
        </g>
        <g
           id="g10022">
          <path
             d="m 1569,1480 h 36 v 0 z m 36,0 v 0 h -36 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10024" />
        </g>
        <g
           id="g10026">
          <path
             d="m 1605,1480 h -36 l 35,-4 z m -36,0 35,-4 h -48 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10028" />
        </g>
        <g
           id="g10030">
          <path
             d="m 1604,1476 h -48 l 48,-6 z m -48,0 48,-6 h -49 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10032" />
        </g>
        <g
           id="g10034">
          <path
             d="m 1580,1470 h -13 l 1,-98 z m -13,0 1,-98 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10036" />
        </g>
        <g
           id="g10038">
          <path
             d="m 1568,1372 h -13 l 12,-5 z m -13,0 12,-5 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10040" />
        </g>
        <g
           id="g10042">
          <path
             d="m 1567,1367 h -13 l 13,-3 z m -13,0 13,-3 h -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10044" />
        </g>
        <g
           id="g10046">
          <path
             d="m 1567,1364 h -13 l 11,-7 z m -13,0 11,-7 h -12 z m 11,-7 h -12 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10048" />
        </g>
        <g
           id="g10050">
          <path
             d="m 1553,1357 h 12 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10052" />
        </g>
        <g
           id="g10054">
          <path
             d="m 1565,1357 h -13 l 10,-7 z m -13,0 10,-7 h -12 z m 10,-7 h -12 z m -12,0 h 12 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10056" />
        </g>
        <g
           id="g10058">
          <path
             d="m 1527,1346 3,-1 h -3 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10060" />
        </g>
        <g
           id="g10062">
          <path
             d="m 1562,1350 h -12 l 9,-5 z m -12,0 9,-5 h -13 z m 9,-5 h -13 z m -13,0 h 13 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10064" />
        </g>
        <g
           id="g10066">
          <path
             d="m 1530,1345 h -3 l 7,-1 z m -3,0 7,-1 h -7 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10068" />
        </g>
        <g
           id="g10070">
          <path
             d="m 1559,1345 h -13 l 12,-2 z m -13,0 12,-2 h -15 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10072" />
        </g>
        <g
           id="g10074">
          <path
             d="m 1534,1344 h -7 l 9,-1 z m -7,0 9,-1 h -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10076" />
        </g>
        <g
           id="g10078">
          <path
             d="m 1558,1343 h -15 14 z m -15,0 h 14 -18 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10080" />
        </g>
        <g
           id="g10082">
          <path
             d="m 1536,1343 h -9 12 z m -9,0 h 12 -13 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10084" />
        </g>
        <g
           id="g10086">
          <path
             d="m 1557,1343 h -31 l 30,-2 z m -31,0 30,-2 h -30 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10088" />
        </g>
        <g
           id="g10090">
          <path
             d="m 1556,1341 h -30 l 25,-4 z m -30,0 25,-4 h -27 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10092" />
        </g>
        <g
           id="g10094">
          <path
             d="m 1551,1337 h -27 l 25,-1 z m -27,0 25,-1 h -25 z m 25,-1 h -25 z m -25,0 h 25 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10096" />
        </g>
        <g
           id="g10098">
          <path
             d="m 1549,1336 h -25 l 23,-1 z m -25,0 23,-1 h -23 z m 23,-1 h -23 z m -23,0 h 23 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10100" />
        </g>
        <g
           id="g10102">
          <path
             d="m 1547,1335 h -23 l 18,-1 z m -23,0 18,-1 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10104" />
        </g>
        <g
           id="g10106">
          <path
             d="m 1530,1334 5,-1 h 6 z m 5,-1 h 6 -5 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10108" />
        </g>
        <g
           id="g10110">
          <path
             d="m 1530,1334 h 12 l -1,-1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10112" />
        </g>
        <path
           d="m 1939,1039 v 0"
           style="fill:none;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path10114" />
        <path
           d="m 1939,1174 v 0"
           style="fill:none;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path10116" />
        <g
           id="g10118">
          <path
             d="m 794,1261 5,-1 h -21 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10120" />
        </g>
        <g
           id="g10122">
          <path
             d="m 799,1260 h -21 l 32,-2 z m -21,0 32,-2 h -39 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10124" />
        </g>
        <g
           id="g10126">
          <path
             d="m 810,1258 h -39 l 45,-2 z m -39,0 45,-2 h -53 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10128" />
        </g>
        <g
           id="g10130">
          <path
             d="m 816,1256 h -53 l 62,-3 z m -53,0 62,-3 h -70 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10132" />
        </g>
        <g
           id="g10134">
          <path
             d="m 825,1253 h -70 l 75,-3 z m -70,0 75,-3 h -82 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10136" />
        </g>
        <g
           id="g10138">
          <path
             d="m 830,1250 h -82 l 91,-5 z m -82,0 91,-5 h -98 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10140" />
        </g>
        <g
           id="g10142">
          <path
             d="m 839,1245 h -98 l 103,-4 z m -98,0 103,-4 H 735 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10144" />
        </g>
        <g
           id="g10146">
          <path
             d="M 844,1241 H 735 l 116,-6 z m -109,0 116,-6 H 729 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10148" />
        </g>
        <g
           id="g10150">
          <path
             d="M 851,1235 H 729 l 126,-5 z m -122,0 126,-5 H 724 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10152" />
        </g>
        <g
           id="g10154">
          <path
             d="M 855,1230 H 724 l 137,-7 z m -131,0 137,-7 H 719 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10156" />
        </g>
        <g
           id="g10158">
          <path
             d="M 861,1223 H 719 l 133,-7 z m -142,0 133,-7 H 715 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10160" />
        </g>
        <g
           id="g10162">
          <path
             d="M 852,1216 H 715 l 135,-2 z m -137,0 135,-2 H 714 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10164" />
        </g>
        <g
           id="g10166">
          <path
             d="m 850,1214 h -62 61 z m -62,0 h 61 -55 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10168" />
        </g>
        <g
           id="g10170">
          <path
             d="m 782,1214 v 0 h -68 z m 0,0 h -68 74 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10172" />
        </g>
        <g
           id="g10174">
          <path
             d="m 849,1214 h -55 l 54,-1 z m -55,0 54,-1 h -48 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10176" />
        </g>
        <g
           id="g10178">
          <path
             d="m 782,1214 h -68 l 63,-2 z m -68,0 63,-2 h -64 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10180" />
        </g>
        <g
           id="g10182">
          <path
             d="m 848,1213 h -48 l 44,-3 z m -48,0 44,-3 h -39 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10184" />
        </g>
        <g
           id="g10186">
          <path
             d="m 777,1212 h -64 l 58,-4 z m -64,0 58,-4 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10188" />
        </g>
        <g
           id="g10190">
          <path
             d="m 844,1210 h -39 l 35,-3 z m -39,0 35,-3 h -30 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10192" />
        </g>
        <g
           id="g10194">
          <path
             d="m 771,1208 h -59 l 55,-3 z m -59,0 55,-3 h -57 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10196" />
        </g>
        <g
           id="g10198">
          <path
             d="m 840,1207 h -30 l 24,-4 z m -30,0 24,-4 h -20 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10200" />
        </g>
        <g
           id="g10202">
          <path
             d="m 767,1205 h -57 l 55,-3 z m -57,0 55,-3 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10204" />
        </g>
        <g
           id="g10206">
          <path
             d="m 765,1202 h -56 l 54,-2 z m -56,0 54,-2 h -55 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10208" />
        </g>
        <g
           id="g10210">
          <path
             d="m 834,1203 h -20 l 13,-5 z m -20,0 13,-5 h -10 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10212" />
        </g>
        <g
           id="g10214">
          <path
             d="m 817,1198 2,-4 h 4 z m 2,-4 h 4 l -3,-2 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10216" />
        </g>
        <g
           id="g10218">
          <path
             d="m 817,1198 h 10 l -4,-4 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10220" />
        </g>
        <g
           id="g10222">
          <path
             d="m 763,1200 h -55 l 53,-6 z m -55,0 53,-6 h -54 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10224" />
        </g>
        <g
           id="g10226">
          <path
             d="m 761,1194 h -54 l 52,-5 z m -54,0 52,-5 h -53 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10228" />
        </g>
        <g
           id="g10230">
          <path
             d="m 759,1189 h -53 l 53,-3 z m -53,0 53,-3 h -54 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10232" />
        </g>
        <g
           id="g10234">
          <path
             d="m 759,1186 h -54 l 54,-3 z m -54,0 54,-3 h -54 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10236" />
        </g>
        <g
           id="g10238">
          <path
             d="m 759,1183 h -54 l 55,-6 z m -54,0 55,-6 h -55 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10240" />
        </g>
        <g
           id="g10242">
          <path
             d="m 760,1177 h -55 l 56,-6 z m -55,0 56,-6 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10244" />
        </g>
        <g
           id="g10246">
          <path
             d="m 761,1171 h -56 l 57,-1 z m -56,0 57,-1 h -57 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10248" />
        </g>
        <g
           id="g10250">
          <path
             d="m 762,1170 h -57 l 59,-4 z m -57,0 59,-4 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10252" />
        </g>
        <g
           id="g10254">
          <path
             d="m 764,1166 h -59 l 63,-5 z m -59,0 63,-5 h -62 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10256" />
        </g>
        <g
           id="g10258">
          <path
             d="m 768,1161 h -62 l 67,-3 z m -62,0 67,-3 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10260" />
        </g>
        <g
           id="g10262">
          <path
             d="m 773,1158 h -66 l 71,-3 z m -66,0 71,-3 h -71 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10264" />
        </g>
        <g
           id="g10266">
          <path
             d="m 779,1155 v 0 h -72 z m 0,0 h -72 71 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10268" />
        </g>
        <g
           id="g10270">
          <path
             d="m 779,1155 h -72 l 77,-2 z m -72,0 77,-2 h -76 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10272" />
        </g>
        <g
           id="g10274">
          <path
             d="m 790,1153 v 0 h -82 z m 0,0 h -82 76 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10276" />
        </g>
        <g
           id="g10278">
          <path
             d="m 790,1153 h -82 l 101,-2 z m -82,0 101,-2 H 709 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10280" />
        </g>
        <g
           id="g10282">
          <path
             d="M 809,1151 H 709 l 118,-6 z m -100,0 118,-6 H 711 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10284" />
        </g>
        <g
           id="g10286">
          <path
             d="M 827,1145 H 711 l 127,-5 z m -116,0 127,-5 H 713 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10288" />
        </g>
        <g
           id="g10290">
          <path
             d="M 838,1140 H 713 l 131,-3 z m -125,0 131,-3 H 714 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10292" />
        </g>
        <g
           id="g10294">
          <path
             d="M 844,1137 H 714 l 144,-11 z m -130,0 144,-11 H 721 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10296" />
        </g>
        <g
           id="g10298">
          <path
             d="M 858,1126 H 721 l 138,-1 z m -137,0 138,-1 H 722 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10300" />
        </g>
        <g
           id="g10302">
          <path
             d="M 859,1125 H 722 l 147,-11 z m -137,0 147,-11 H 731 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10304" />
        </g>
        <g
           id="g10306">
          <path
             d="M 869,1114 H 731 l 141,-3 z m -138,0 141,-3 H 736 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10308" />
        </g>
        <g
           id="g10310">
          <path
             d="M 872,1111 H 736 l 139,-7 z m -136,0 139,-7 H 744 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10312" />
        </g>
        <g
           id="g10314">
          <path
             d="M 875,1104 H 744 l 135,-7 z m -131,0 135,-7 H 758 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10316" />
        </g>
        <g
           id="g10318">
          <path
             d="M 879,1097 H 758 l 123,-3 z m -121,0 123,-3 H 768 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10320" />
        </g>
        <g
           id="g10322">
          <path
             d="M 881,1094 H 768 l 114,-2 z m -113,0 114,-2 H 773 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10324" />
        </g>
        <g
           id="g10326">
          <path
             d="M 882,1092 H 773 l 109,-1 z m -109,0 109,-1 h -93 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10328" />
        </g>
        <g
           id="g10330">
          <path
             d="m 882,1091 h -93 l 93,-1 z m -93,0 93,-1 h -86 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10332" />
        </g>
        <g
           id="g10334">
          <path
             d="m 882,1090 h -86 l 87,-2 z m -86,0 87,-2 h -80 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10336" />
        </g>
        <g
           id="g10338">
          <path
             d="m 883,1088 h -80 l 81,-3 z m -80,0 81,-3 h -74 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10340" />
        </g>
        <g
           id="g10342">
          <path
             d="m 884,1085 h -74 l 76,-4 z m -74,0 76,-4 h -70 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10344" />
        </g>
        <g
           id="g10346">
          <path
             d="m 886,1081 h -70 l 71,-5 z m -70,0 71,-5 h -67 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10348" />
        </g>
        <g
           id="g10350">
          <path
             d="m 887,1076 h -67 l 68,-1 z m -67,0 68,-1 h -67 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10352" />
        </g>
        <g
           id="g10354">
          <path
             d="m 888,1075 h -67 l 67,-6 z m -67,0 67,-6 h -63 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10356" />
        </g>
        <g
           id="g10358">
          <path
             d="m 888,1069 h -63 l 64,-7 z m -63,0 64,-7 h -62 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10360" />
        </g>
        <g
           id="g10362">
          <path
             d="m 889,1062 h -62 l 63,-5 z m -62,0 63,-5 h -62 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10364" />
        </g>
        <g
           id="g10366">
          <path
             d="m 890,1057 h -62 l 62,-2 z m -62,0 62,-2 h -62 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10368" />
        </g>
        <g
           id="g10370">
          <path
             d="m 890,1055 h -62 l 62,-7 z m -62,0 62,-7 h -62 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10372" />
        </g>
        <g
           id="g10374">
          <path
             d="m 890,1048 h -62 l 61,-7 z m -62,0 61,-7 h -62 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10376" />
        </g>
        <g
           id="g10378">
          <path
             d="m 889,1041 h -62 l 62,-3 z m -62,0 62,-3 h -63 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10380" />
        </g>
        <g
           id="g10382">
          <path
             d="m 754,1038 2,-4 h -8 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10384" />
        </g>
        <g
           id="g10386">
          <path
             d="m 889,1038 h -63 l 62,-4 z m -63,0 62,-4 h -64 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10388" />
        </g>
        <g
           id="g10390">
          <path
             d="m 756,1034 h -8 l 9,-3 z m -8,0 9,-3 h -12 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10392" />
        </g>
        <g
           id="g10394">
          <path
             d="m 888,1034 h -64 l 63,-6 z m -64,0 63,-6 h -67 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10396" />
        </g>
        <g
           id="g10398">
          <path
             d="m 757,1031 h -12 l 17,-5 z m -12,0 17,-5 h -25 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10400" />
        </g>
        <g
           id="g10402">
          <path
             d="m 887,1028 h -67 l 66,-5 z m -67,0 66,-5 h -71 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10404" />
        </g>
        <g
           id="g10406">
          <path
             d="m 762,1026 h -25 l 30,-5 z m -25,0 30,-5 h -37 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10408" />
        </g>
        <g
           id="g10410">
          <path
             d="m 886,1023 h -71 l 70,-4 z m -71,0 70,-4 h -75 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10412" />
        </g>
        <g
           id="g10414">
          <path
             d="m 885,1019 h -75 l 74,-1 z m -75,0 74,-1 h -75 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10416" />
        </g>
        <g
           id="g10418">
          <path
             d="m 767,1021 h -37 l 43,-4 z m -37,0 43,-4 h -48 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10420" />
        </g>
        <g
           id="g10422">
          <path
             d="m 884,1018 h -75 l 74,-3 z m -75,0 74,-3 h -81 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10424" />
        </g>
        <g
           id="g10426">
          <path
             d="m 773,1017 h -48 l 55,-2 z m -48,0 55,-2 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10428" />
        </g>
        <g
           id="g10430">
          <path
             d="m 883,1015 h -81 l 80,-1 z m -81,0 80,-1 h -87 z m 80,-1 h -87 -7 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10432" />
        </g>
        <g
           id="g10434">
          <path
             d="m 795,1014 h 87 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10436" />
        </g>
        <g
           id="g10438">
          <path
             d="m 780,1015 h -59 l 67,-1 z m -59,0 67,-1 h -68 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10440" />
        </g>
        <g
           id="g10442">
          <path
             d="M 882,1014 H 720 l 157,-12 z m -162,0 157,-12 H 704 Z m 157,-12 h -173 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10444" />
        </g>
        <g
           id="g10446">
          <path
             d="m 704,1002 h 173 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10448" />
        </g>
        <g
           id="g10450">
          <path
             d="M 877,1002 H 703 l 163,-16 z m -174,0 163,-16 H 714 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10452" />
        </g>
        <g
           id="g10454">
          <path
             d="m 865,986 v 0 H 714 Z m 0,0 H 714 866 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10456" />
        </g>
        <g
           id="g10458">
          <path
             d="M 865,986 H 714 l 138,-13 z m -151,0 138,-13 H 728 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10460" />
        </g>
        <g
           id="g10462">
          <path
             d="m 851,973 v 0 H 728 Z m 0,0 H 728 852 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10464" />
        </g>
        <g
           id="g10466">
          <path
             d="M 851,973 H 728 l 108,-10 z m -123,0 108,-10 h -92 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10468" />
        </g>
        <g
           id="g10470">
          <path
             d="m 835,963 v 0 h -91 z m 0,0 h -91 92 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10472" />
        </g>
        <g
           id="g10474">
          <path
             d="m 835,963 h -91 l 74,-7 z m -91,0 74,-7 h -57 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10476" />
        </g>
        <g
           id="g10478">
          <path
             d="m 818,956 h -57 56 z m -57,0 h 56 -55 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10480" />
        </g>
        <g
           id="g10482">
          <path
             d="m 762,956 18,-4 h 20 z m 18,-4 h 20 -19 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10484" />
        </g>
        <g
           id="g10486">
          <path
             d="m 762,956 h 55 l -17,-4 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10488" />
        </g>
        <g
           id="g10490">
          <path
             d="m 1287,1261 149,-122 h -149 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10492" />
        </g>
        <g
           id="g10494">
          <path
             d="m 1427,1074 h 149 V 952 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10496" />
        </g>
        <g
           id="g10498">
          <path
             d="m 1576,1261 h -61 l 61,-187 z m -61,0 61,-187 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10500" />
        </g>
        <g
           id="g10502">
          <path
             d="m 1436,1139 h -88 l 167,-65 z m -88,0 167,-65 h -88 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10504" />
        </g>
        <g
           id="g10506">
          <path
             d="m 1348,1139 h -61 l 61,-65 z m -61,0 61,-65 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10508" />
        </g>
        <g
           id="g10510">
          <path
             d="m 1348,1074 h -61 l 61,-122 z m -61,0 61,-122 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10512" />
        </g>
        <g
           id="g10514">
          <path
             d="m 2076,1261 h 65 l -65,-309 z m 65,0 -65,-309 h 65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10516" />
        </g>
        <g
           id="g10518">
          <path
             d="m 2371,1261 h -157 l 157,-60 z m -157,0 157,-60 h -157 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10520" />
        </g>
        <g
           id="g10522">
          <path
             d="m 2275,1201 h -61 l 61,-60 z m -61,0 61,-60 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10524" />
        </g>
        <g
           id="g10526">
          <path
             d="m 2385,1141 h -171 l 171,-59 z m -171,0 171,-59 h -171 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10528" />
        </g>
        <g
           id="g10530">
          <path
             d="m 2275,1082 h -61 l 61,-71 z m -61,0 61,-71 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10532" />
        </g>
        <g
           id="g10534">
          <path
             d="m 2405,1011 h -191 l 191,-59 z m -191,0 191,-59 h -191 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10536" />
        </g>
        <g
           id="g10538">
          <path
             d="m 2593,1261 h 4 -6 z m 4,0 h -6 -4 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10540" />
        </g>
        <g
           id="g10542">
          <path
             d="m 2591,1261 h 6 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10544" />
        </g>
        <g
           id="g10546">
          <path
             d="m 2597,1261 h -10 l 20,-1 z m -10,0 20,-1 h -30 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10548" />
        </g>
        <g
           id="g10550">
          <path
             d="m 2607,1260 h -30 34 z m -30,0 h 34 -36 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10552" />
        </g>
        <g
           id="g10554">
          <path
             d="m 2611,1260 h -36 l 49,-2 z m -36,0 49,-2 h -63 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10556" />
        </g>
        <g
           id="g10558">
          <path
             d="m 2624,1258 h -63 65 z m -63,0 h 65 -69 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10560" />
        </g>
        <g
           id="g10562">
          <path
             d="m 2626,1258 h -69 l 80,-3 z m -69,0 80,-3 h -90 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10564" />
        </g>
        <g
           id="g10566">
          <path
             d="m 2637,1255 h -90 l 96,-2 z m -90,0 96,-2 h -105 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10568" />
        </g>
        <g
           id="g10570">
          <path
             d="m 2643,1253 h -105 l 111,-2 z m -105,0 111,-2 h -116 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10572" />
        </g>
        <g
           id="g10574">
          <path
             d="m 2649,1251 h -116 l 127,-4 z m -116,0 127,-4 h -139 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10576" />
        </g>
        <g
           id="g10578">
          <path
             d="m 2660,1247 h -139 l 139,-1 z m -139,0 139,-1 h -140 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10580" />
        </g>
        <g
           id="g10582">
          <path
             d="m 2660,1246 h -140 l 151,-6 z m -140,0 151,-6 h -162 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10584" />
        </g>
        <g
           id="g10586">
          <path
             d="m 2671,1240 h -162 l 165,-2 z m -162,0 165,-2 h -169 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10588" />
        </g>
        <g
           id="g10590">
          <path
             d="m 2674,1238 h -169 l 176,-4 z m -169,0 176,-4 h -183 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10592" />
        </g>
        <g
           id="g10594">
          <path
             d="m 2681,1234 h -183 l 190,-6 z m -183,0 190,-6 h -197 z m 190,-6 h -197 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10596" />
        </g>
        <g
           id="g10598">
          <path
             d="m 2491,1228 h 197 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10600" />
        </g>
        <g
           id="g10602">
          <path
             d="m 2688,1228 h -198 l 210,-12 z m -198,0 210,-12 h -223 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10604" />
        </g>
        <g
           id="g10606">
          <path
             d="m 2700,1216 h -223 l 224,-2 z m -223,0 224,-2 h -225 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10608" />
        </g>
        <g
           id="g10610">
          <path
             d="m 2701,1214 h -225 l 227,-1 z m -225,0 227,-1 h -229 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10612" />
        </g>
        <g
           id="g10614">
          <path
             d="m 2590,1213 h 113 v 0 z m 113,0 v 0 h -113 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10616" />
        </g>
        <g
           id="g10618">
          <path
             d="m 2474,1213 h 116 v 0 z m 116,0 v 0 h -116 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10620" />
        </g>
        <g
           id="g10622">
          <path
             d="m 2590,1213 h -116 l 101,-1 z m -116,0 101,-1 h -102 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10624" />
        </g>
        <g
           id="g10626">
          <path
             d="m 2703,1213 h -113 l 114,-2 z m -113,0 114,-2 h -100 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10628" />
        </g>
        <g
           id="g10630">
          <path
             d="m 2575,1212 h -102 l 92,-3 z m -102,0 92,-3 h -93 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10632" />
        </g>
        <g
           id="g10634">
          <path
             d="m 2565,1209 h -93 90 z m -93,0 h 90 -91 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10636" />
        </g>
        <g
           id="g10638">
          <path
             d="m 2704,1211 h -100 l 102,-3 z m -100,0 102,-3 h -88 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10640" />
        </g>
        <g
           id="g10642">
          <path
             d="m 2562,1209 h -91 l 78,-6 z m -91,0 78,-6 h -82 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10644" />
        </g>
        <g
           id="g10646">
          <path
             d="m 2549,1203 h -82 81 z m -82,0 h 81 -82 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10648" />
        </g>
        <g
           id="g10650">
          <path
             d="m 2706,1208 h -88 l 92,-6 z m -88,0 92,-6 h -79 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10652" />
        </g>
        <g
           id="g10654">
          <path
             d="m 2710,1202 h -79 l 82,-4 z m -79,0 82,-4 h -76 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10656" />
        </g>
        <g
           id="g10658">
          <path
             d="m 2548,1203 h -82 l 71,-7 z m -82,0 71,-7 h -75 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10660" />
        </g>
        <g
           id="g10662">
          <path
             d="m 2713,1198 h -76 l 79,-4 z m -76,0 79,-4 h -73 z m 79,-4 h -73 z m -73,0 h 73 v 0 z m 73,0 v 0 h -73 z m 0,0 h -73 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10664" />
        </g>
        <g
           id="g10666">
          <path
             d="m 2537,1196 h -75 l 68,-6 z m -75,0 68,-6 h -72 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10668" />
        </g>
        <g
           id="g10670">
          <path
             d="m 2530,1190 h -72 l 69,-3 z m -72,0 69,-3 h -71 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10672" />
        </g>
        <g
           id="g10674">
          <path
             d="m 2716,1194 h -73 l 77,-8 z m -73,0 77,-8 h -69 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10676" />
        </g>
        <g
           id="g10678">
          <path
             d="m 2720,1186 h -69 l 73,-7 z m -69,0 73,-7 h -67 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10680" />
        </g>
        <g
           id="g10682">
          <path
             d="m 2724,1179 h -67 l 65,-1 z m -67,0 65,-1 h -64 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10684" />
        </g>
        <g
           id="g10686">
          <path
             d="m 2527,1187 h -71 l 62,-11 z m -71,0 62,-11 h -68 z m 62,-11 h -68 z m -68,0 h 68 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10688" />
        </g>
        <g
           id="g10690">
          <path
             d="m 2722,1178 h -64 l 39,-10 z m -64,0 39,-10 h -33 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10692" />
        </g>
        <g
           id="g10694">
          <path
             d="m 2518,1176 h -68 l 60,-12 z m -68,0 60,-12 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10696" />
        </g>
        <g
           id="g10698">
          <path
             d="m 2664,1168 3,-7 h 14 z m 3,-7 h 14 l -12,-4 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10700" />
        </g>
        <g
           id="g10702">
          <path
             d="m 2664,1168 h 33 l -16,-7 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10704" />
        </g>
        <g
           id="g10706">
          <path
             d="m 2510,1164 h -65 l 64,-3 z m -65,0 64,-3 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10708" />
        </g>
        <g
           id="g10710">
          <path
             d="m 2509,1161 h -65 l 60,-11 z m -65,0 60,-11 h -63 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10712" />
        </g>
        <g
           id="g10714">
          <path
             d="m 2504,1150 h -63 l 62,-4 z m -63,0 62,-4 h -63 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10716" />
        </g>
        <g
           id="g10718">
          <path
             d="m 2503,1146 h -63 l 60,-7 z m -63,0 60,-7 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10720" />
        </g>
        <g
           id="g10722">
          <path
             d="m 2500,1139 h -61 l 59,-9 z m -61,0 59,-9 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10724" />
        </g>
        <g
           id="g10726">
          <path
             d="m 2498,1130 h -61 l 61,-2 z m -61,0 61,-2 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10728" />
        </g>
        <g
           id="g10730">
          <path
             d="m 2498,1128 h -61 l 59,-12 z m -61,0 59,-12 h -60 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10732" />
        </g>
        <g
           id="g10734">
          <path
             d="m 2496,1116 h -60 l 60,-3 z m -60,0 60,-3 h -60 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10736" />
        </g>
        <g
           id="g10738">
          <path
             d="m 2496,1113 h -60 l 60,-8 z m -60,0 60,-8 h -60 z m 60,-8 h -60 z m -60,0 h 60 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10740" />
        </g>
        <g
           id="g10742">
          <path
             d="m 2740,1122 h -150 l 149,-25 z m -150,0 149,-25 h -149 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10744" />
        </g>
        <g
           id="g10746">
          <path
             d="m 2496,1105 h -60 l 60,-9 z m -60,0 60,-9 h -60 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10748" />
        </g>
        <g
           id="g10750">
          <path
             d="m 2496,1096 h -60 l 60,-3 z m -60,0 60,-3 h -60 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10752" />
        </g>
        <g
           id="g10754">
          <path
             d="m 2496,1093 h -60 l 62,-11 z m -60,0 62,-11 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10756" />
        </g>
        <g
           id="g10758">
          <path
             d="m 2498,1082 h -61 l 61,-2 z m -61,0 61,-2 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10760" />
        </g>
        <g
           id="g10762">
          <path
             d="m 2739,1097 h -149 l 146,-23 z m -149,0 146,-23 h -146 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10764" />
        </g>
        <g
           id="g10766">
          <path
             d="m 2736,1074 h -146 l 146,-2 z m -146,0 146,-2 h -146 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10768" />
        </g>
        <g
           id="g10770">
          <path
             d="m 2498,1080 h -61 l 63,-9 z m -61,0 63,-9 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10772" />
        </g>
        <g
           id="g10774">
          <path
             d="m 2500,1071 h -61 l 63,-5 z m -61,0 63,-5 h -62 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10776" />
        </g>
        <g
           id="g10778">
          <path
             d="m 2502,1066 h -62 l 63,-6 z m -62,0 63,-6 h -62 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10780" />
        </g>
        <g
           id="g10782">
          <path
             d="m 2736,1072 h -58 l 55,-15 z m -58,0 55,-15 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10784" />
        </g>
        <g
           id="g10786">
          <path
             d="m 2733,1057 h -59 l 58,-3 z m -59,0 58,-3 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10788" />
        </g>
        <g
           id="g10790">
          <path
             d="m 2503,1060 h -62 l 66,-9 z m -62,0 66,-9 h -64 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10792" />
        </g>
        <g
           id="g10794">
          <path
             d="m 2507,1051 h -64 l 65,-1 z m -64,0 65,-1 h -64 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10796" />
        </g>
        <g
           id="g10798">
          <path
             d="m 2732,1054 h -59 l 56,-8 z m -59,0 56,-8 h -60 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10800" />
        </g>
        <g
           id="g10802">
          <path
             d="m 2729,1046 h -60 l 59,-3 z m -60,0 59,-3 h -60 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10804" />
        </g>
        <g
           id="g10806">
          <path
             d="m 2508,1050 h -64 l 69,-9 z m -64,0 69,-9 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10808" />
        </g>
        <g
           id="g10810">
          <path
             d="m 2513,1041 h -65 l 67,-3 z m -65,0 67,-3 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10812" />
        </g>
        <g
           id="g10814">
          <path
             d="m 2728,1043 h -60 l 57,-9 z m -60,0 57,-9 h -63 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10816" />
        </g>
        <g
           id="g10818">
          <path
             d="m 2515,1038 h -66 l 71,-6 z m -66,0 71,-6 h -68 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10820" />
        </g>
        <g
           id="g10822">
          <path
             d="m 2725,1034 h -63 l 61,-4 z m -63,0 61,-4 h -63 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10824" />
        </g>
        <g
           id="g10826">
          <path
             d="m 2520,1032 h -68 l 73,-7 z m -68,0 73,-7 h -70 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10828" />
        </g>
        <g
           id="g10830">
          <path
             d="m 2525,1025 h -70 l 72,-2 z m -70,0 72,-2 h -71 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10832" />
        </g>
        <g
           id="g10834">
          <path
             d="m 2723,1030 h -63 l 59,-8 z m -63,0 59,-8 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10836" />
        </g>
        <g
           id="g10838">
          <path
             d="m 2650,1019 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10840" />
        </g>
        <g
           id="g10842">
          <path
             d="m 2719,1022 h -66 l 64,-3 z m -66,0 64,-3 h -67 z m 64,-3 h -67 z m -67,0 h 67 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10844" />
        </g>
        <g
           id="g10846">
          <path
             d="m 2527,1023 h -71 l 83,-10 z m -71,0 83,-10 h -76 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10848" />
        </g>
        <g
           id="g10850">
          <path
             d="m 2539,1013 h -76 l 77,-1 z m -76,0 77,-1 h -76 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10852" />
        </g>
        <g
           id="g10854">
          <path
             d="m 2717,1019 h -67 l 62,-8 z m -67,0 62,-8 h -71 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10856" />
        </g>
        <g
           id="g10858">
          <path
             d="m 2712,1011 h -71 l 70,-2 z m -71,0 70,-2 h -73 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10860" />
        </g>
        <g
           id="g10862">
          <path
             d="m 2540,1012 h -76 l 85,-5 z m -76,0 85,-5 h -82 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10864" />
        </g>
        <g
           id="g10866">
          <path
             d="m 2549,1007 h -82 l 89,-4 z m -82,0 89,-4 h -86 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10868" />
        </g>
        <g
           id="g10870">
          <path
             d="m 2711,1009 h -73 l 68,-7 z m -73,0 68,-7 h -82 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10872" />
        </g>
        <g
           id="g10874">
          <path
             d="m 2706,1002 h -82 l 81,-1 z m -82,0 81,-1 h -83 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10876" />
        </g>
        <g
           id="g10878">
          <path
             d="m 2556,1003 h -86 l 99,-3 z m -86,0 99,-3 h -96 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10880" />
        </g>
        <g
           id="g10882">
          <path
             d="m 2569,1000 h -96 l 100,-2 z m -96,0 100,-2 h -99 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10884" />
        </g>
        <g
           id="g10886">
          <path
             d="m 2705,1001 h -83 l 80,-3 z m -83,0 80,-3 h -94 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10888" />
        </g>
        <g
           id="g10890">
          <path
             d="m 2702,998 h -94 l 93,-1 z m -94,0 93,-1 h -109 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10892" />
        </g>
        <g
           id="g10894">
          <path
             d="m 2573,998 h -99 l 118,-1 z m -99,0 118,-1 h -116 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10896" />
        </g>
        <g
           id="g10898">
          <path
             d="m 2701,997 h -225 l 221,-5 z m -225,0 221,-5 h -217 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10900" />
        </g>
        <g
           id="g10902">
          <path
             d="m 2697,992 h -217 l 210,-6 z m -217,0 210,-6 h -203 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10904" />
        </g>
        <g
           id="g10906">
          <path
             d="m 2690,986 h -203 l 201,-2 z m -203,0 201,-2 h -198 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10908" />
        </g>
        <g
           id="g10910">
          <path
             d="m 2688,984 h -198 l 188,-7 z m -198,0 188,-7 h -178 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10912" />
        </g>
        <g
           id="g10914">
          <path
             d="m 2678,977 h -178 l 176,-2 z m -178,0 176,-2 h -174 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10916" />
        </g>
        <g
           id="g10918">
          <path
             d="m 2676,975 h -174 l 166,-5 z m -174,0 166,-5 h -157 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10920" />
        </g>
        <g
           id="g10922">
          <path
             d="m 2668,970 h -157 l 149,-4 z m -157,0 149,-4 h -142 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10924" />
        </g>
        <g
           id="g10926">
          <path
             d="m 2660,966 h -142 l 139,-1 z m -142,0 139,-1 h -136 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10928" />
        </g>
        <g
           id="g10930">
          <path
             d="m 2657,965 h -136 l 125,-5 z m -136,0 125,-5 h -113 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10932" />
        </g>
        <g
           id="g10934">
          <path
             d="m 2646,960 h -113 l 109,-1 z m -113,0 109,-1 h -106 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10936" />
        </g>
        <g
           id="g10938">
          <path
             d="m 2642,959 h -106 l 98,-2 z m -106,0 98,-2 h -88 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10940" />
        </g>
        <g
           id="g10942">
          <path
             d="m 2634,957 h -88 l 78,-2 z m -88,0 78,-2 h -69 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10944" />
        </g>
        <g
           id="g10946">
          <path
             d="m 2624,955 h -69 l 66,-1 z m -69,0 66,-1 h -62 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10948" />
        </g>
        <g
           id="g10950">
          <path
             d="m 2621,954 h -62 l 50,-2 z m -62,0 50,-2 h -36 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10952" />
        </g>
        <g
           id="g10954">
          <path
             d="m 2609,952 h -36 30 z m -36,0 h 30 -27 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10956" />
        </g>
        <g
           id="g10958">
          <path
             d="m 2603,952 h -27 19 z m -27,0 h 19 -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10960" />
        </g>
        <g
           id="g10962">
          <path
             d="m 2586,952 h 1 7 z m 1,0 h 7 -2 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10964" />
        </g>
        <g
           id="g10966">
          <path
             d="m 2586,952 h 9 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10968" />
        </g>
        <path
           d="m 1136,1047 28,-53"
           style="fill:none;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path10970" />
        <g
           id="g10972">
          <path
             d="m 1090,1261 65,-124 h -130 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10974" />
        </g>
        <g
           id="g10976">
          <path
             d="m 1155,1137 h -66 l 112,-90 z m -66,0 112,-90 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10978" />
        </g>
        <g
           id="g10980">
          <path
             d="m 1089,1137 h -64 l 17,-90 z m -64,0 17,-90 h -64 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10982" />
        </g>
        <g
           id="g10984">
          <path
             d="m 1201,1047 h -65 l 93,-53 z m -65,0 93,-53 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10986" />
        </g>
        <g
           id="g10988">
          <path
             d="M 1136,1047 H 978 l 186,-53 z m -158,0 186,-53 H 950 Z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10990" />
        </g>
        <g
           id="g10992">
          <path
             d="m 1229,994 h -65 l 87,-42 z m -65,0 87,-42 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10994" />
        </g>
        <g
           id="g10996">
          <path
             d="m 1014,994 h -64 l 42,-42 z m -64,0 42,-42 h -64 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path10998" />
        </g>
        <g
           id="g11000">
          <path
             d="m 1872,1261 h -126 l 143,-1 z m -126,0 143,-1 h -143 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11002" />
        </g>
        <g
           id="g11004">
          <path
             d="m 1889,1260 h -143 l 158,-3 z m -143,0 158,-3 h -158 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11006" />
        </g>
        <g
           id="g11008">
          <path
             d="m 1904,1257 h -158 l 173,-4 z m -158,0 173,-4 h -173 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11010" />
        </g>
        <g
           id="g11012">
          <path
             d="m 1919,1253 h -173 l 188,-6 z m -173,0 188,-6 h -188 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11014" />
        </g>
        <g
           id="g11016">
          <path
             d="m 1934,1247 h -188 l 202,-7 z m -188,0 202,-7 h -202 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11018" />
        </g>
        <g
           id="g11020">
          <path
             d="m 1948,1240 h -202 l 216,-9 z m -202,0 216,-9 h -216 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11022" />
        </g>
        <g
           id="g11024">
          <path
             d="m 1962,1231 h -216 l 228,-11 z m -216,0 228,-11 h -228 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11026" />
        </g>
        <g
           id="g11028">
          <path
             d="m 1974,1220 h -228 l 235,-7 z m -228,0 235,-7 h -235 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11030" />
        </g>
        <g
           id="g11032">
          <path
             d="m 1981,1213 h -128 129 z m -128,0 h 129 -116 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11034" />
        </g>
        <g
           id="g11036">
          <path
             d="m 1982,1213 h -116 l 118,-2 z m -116,0 118,-2 h -106 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11038" />
        </g>
        <g
           id="g11040">
          <path
             d="m 1984,1211 h -106 l 107,-2 z m -106,0 107,-2 h -100 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11042" />
        </g>
        <g
           id="g11044">
          <path
             d="m 1985,1209 h -100 l 101,-1 z m -100,0 101,-1 h -96 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11046" />
        </g>
        <g
           id="g11048">
          <path
             d="m 1986,1208 h -96 l 100,-4 z m -96,0 100,-4 h -88 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11050" />
        </g>
        <g
           id="g11052">
          <path
             d="m 1990,1204 h -88 l 92,-6 z m -88,0 92,-6 h -82 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11054" />
        </g>
        <g
           id="g11056">
          <path
             d="m 1994,1198 h -82 l 83,-1 z m -82,0 83,-1 h -81 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11058" />
        </g>
        <g
           id="g11060">
          <path
             d="m 1995,1197 h -81 l 85,-6 z m -81,0 85,-6 h -77 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11062" />
        </g>
        <g
           id="g11064">
          <path
             d="m 1999,1191 h -77 l 82,-8 z m -77,0 82,-8 h -73 z m 82,-8 h -73 z m -73,0 h 73 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11066" />
        </g>
        <g
           id="g11068">
          <path
             d="m 2004,1183 h -73 l 77,-7 z m -73,0 77,-7 h -71 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11070" />
        </g>
        <g
           id="g11072">
          <path
             d="m 2008,1176 h -71 l 72,-2 z m -71,0 72,-2 h -70 z m 72,-2 h -70 z m -70,0 h 70 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11074" />
        </g>
        <g
           id="g11076">
          <path
             d="m 2009,1174 h -70 l 72,-4 z m -70,0 72,-4 h -69 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11078" />
        </g>
        <g
           id="g11080">
          <path
             d="m 2011,1170 h -69 l 73,-11 z m -69,0 73,-11 h -67 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11082" />
        </g>
        <g
           id="g11084">
          <path
             d="m 2015,1159 h -67 l 68,-2 z m -67,0 68,-2 h -67 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11086" />
        </g>
        <g
           id="g11088">
          <path
             d="m 2016,1157 h -67 l 71,-12 z m -67,0 71,-12 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11090" />
        </g>
        <g
           id="g11092">
          <path
             d="m 2020,1145 h -66 l 66,-3 z m -66,0 66,-3 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11094" />
        </g>
        <g
           id="g11096">
          <path
             d="m 2020,1142 h -65 l 68,-10 z m -65,0 68,-10 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11098" />
        </g>
        <g
           id="g11100">
          <path
             d="m 2023,1132 h -65 l 66,-7 z m -65,0 66,-7 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11102" />
        </g>
        <g
           id="g11104">
          <path
             d="m 2024,1125 h -65 l 65,-6 z m -65,0 65,-6 h -64 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11106" />
        </g>
        <g
           id="g11108">
          <path
             d="m 2024,1119 h -64 l 65,-13 z m -64,0 65,-13 h -64 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11110" />
        </g>
        <g
           id="g11112">
          <path
             d="m 2025,1106 h -64 l 63,-17 z m -64,0 63,-17 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11114" />
        </g>
        <g
           id="g11116">
          <path
             d="m 2024,1089 h -65 l 65,-1 z m -65,0 65,-1 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11118" />
        </g>
        <g
           id="g11120">
          <path
             d="m 2024,1088 h -65 l 62,-17 z m -65,0 62,-17 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11122" />
        </g>
        <g
           id="g11124">
          <path
             d="m 2021,1071 h -66 l 66,-1 z m -66,0 66,-1 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11126" />
        </g>
        <g
           id="g11128">
          <path
             d="m 2021,1070 h -66 l 61,-16 z m -66,0 61,-16 h -67 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11130" />
        </g>
        <g
           id="g11132">
          <path
             d="m 2016,1054 h -67 66 z m -67,0 h 66 -67 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11134" />
        </g>
        <g
           id="g11136">
          <path
             d="m 2015,1054 h -67 l 61,-15 z m -67,0 61,-15 h -70 z m 61,-15 h -70 z m -70,0 h 70 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11138" />
        </g>
        <g
           id="g11140">
          <path
             d="m 2009,1039 h -70 l 69,-1 z m -70,0 69,-1 h -70 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11142" />
        </g>
        <g
           id="g11144">
          <path
             d="m 2008,1038 h -70 l 66,-8 z m -70,0 66,-8 h -73 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11146" />
        </g>
        <g
           id="g11148">
          <path
             d="m 2004,1030 h -73 l 68,-8 z m -73,0 68,-8 h -76 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11150" />
        </g>
        <g
           id="g11152">
          <path
             d="m 1999,1022 h -76 l 76,-1 z m -76,0 76,-1 h -77 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11154" />
        </g>
        <g
           id="g11156">
          <path
             d="m 1999,1021 h -77 l 72,-6 z m -77,0 72,-6 h -82 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11158" />
        </g>
        <g
           id="g11160">
          <path
             d="m 1994,1015 h -82 l 78,-6 z m -82,0 78,-6 h -88 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11162" />
        </g>
        <g
           id="g11164">
          <path
             d="m 1990,1009 h -88 l 86,-2 z m -88,0 86,-2 h -91 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11166" />
        </g>
        <g
           id="g11168">
          <path
             d="m 1988,1007 h -91 l 89,-2 z m -91,0 89,-2 h -96 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11170" />
        </g>
        <g
           id="g11172">
          <path
             d="m 1986,1005 h -96 l 93,-3 z m -96,0 93,-3 h -105 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11174" />
        </g>
        <g
           id="g11176">
          <path
             d="m 1983,1002 h -105 l 104,-2 z m -105,0 104,-2 h -116 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11178" />
        </g>
        <g
           id="g11180">
          <path
             d="m 1807,1213 h -61 l 61,-214 z m -61,0 61,-214 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11182" />
        </g>
        <g
           id="g11184">
          <path
             d="m 1982,1000 h -116 l 115,-1 z m -116,0 115,-1 h -128 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11186" />
        </g>
        <g
           id="g11188">
          <path
             d="m 1981,999 h -235 l 230,-5 z m -235,0 230,-5 h -230 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11190" />
        </g>
        <g
           id="g11192">
          <path
             d="m 1976,994 h -230 l 217,-12 z m -230,0 217,-12 h -217 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11194" />
        </g>
        <g
           id="g11196">
          <path
             d="m 1963,982 h -217 l 202,-10 z m -217,0 202,-10 h -202 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11198" />
        </g>
        <g
           id="g11200">
          <path
             d="m 1948,972 h -202 l 186,-8 z m -202,0 186,-8 h -186 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11202" />
        </g>
        <g
           id="g11204">
          <path
             d="m 1932,964 h -186 l 178,-3 z m -186,0 178,-3 h -178 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11206" />
        </g>
        <g
           id="g11208">
          <path
             d="m 1924,961 h -178 l 175,-1 z m -178,0 175,-1 h -175 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11210" />
        </g>
        <g
           id="g11212">
          <path
             d="m 1921,960 h -175 l 172,-1 z m -175,0 172,-1 h -172 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11214" />
        </g>
        <g
           id="g11216">
          <path
             d="m 1918,959 h -172 l 163,-3 z m -172,0 163,-3 h -163 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11218" />
        </g>
        <g
           id="g11220">
          <path
             d="m 1909,956 h -163 l 145,-3 z m -163,0 145,-3 h -145 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11222" />
        </g>
        <g
           id="g11224">
          <path
             d="m 1891,953 h -145 l 126,-1 z m -145,0 126,-1 h -126 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11226" />
        </g>
        <g
           id="g11228">
          <path
             d="m 2959,1261 24,-2 h -48 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11230" />
        </g>
        <g
           id="g11232">
          <path
             d="m 2983,1259 h -48 l 72,-5 z m -48,0 72,-5 h -96 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11234" />
        </g>
        <g
           id="g11236">
          <path
             d="m 3007,1254 h -96 l 118,-10 z m -96,0 118,-10 h -140 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11238" />
        </g>
        <g
           id="g11240">
          <path
             d="m 3029,1244 h -140 l 161,-12 z m -140,0 161,-12 h -182 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11242" />
        </g>
        <g
           id="g11244">
          <path
             d="m 3050,1232 h -182 l 201,-16 z m -182,0 201,-16 h -219 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11246" />
        </g>
        <g
           id="g11248">
          <path
             d="m 3069,1216 h -219 l 226,-9 z m -219,0 226,-9 h -234 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11250" />
        </g>
        <g
           id="g11252">
          <path
             d="m 3076,1207 h -117 l 119,-2 z m -117,0 119,-2 h -99 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11254" />
        </g>
        <g
           id="g11256">
          <path
             d="m 2959,1207 h -117 l 98,-2 z m -117,0 98,-2 h -99 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11258" />
        </g>
        <g
           id="g11260">
          <path
             d="m 3078,1205 h -99 l 104,-6 z m -99,0 104,-6 h -85 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11262" />
        </g>
        <g
           id="g11264">
          <path
             d="m 2940,1205 h -99 l 80,-6 z m -99,0 80,-6 h -85 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11266" />
        </g>
        <g
           id="g11268">
          <path
             d="m 3083,1199 h -85 l 86,-2 z m -85,0 86,-2 h -83 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11270" />
        </g>
        <g
           id="g11272">
          <path
             d="m 2921,1199 h -85 l 81,-2 z m -85,0 81,-2 h -83 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11274" />
        </g>
        <g
           id="g11276">
          <path
             d="m 3084,1197 h -83 l 88,-7 z m -83,0 88,-7 h -74 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11278" />
        </g>
        <g
           id="g11280">
          <path
             d="m 2917,1197 h -83 l 69,-7 z m -83,0 69,-7 h -73 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11282" />
        </g>
        <g
           id="g11284">
          <path
             d="m 3089,1190 h -74 l 81,-12 z m -74,0 81,-12 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11286" />
        </g>
        <g
           id="g11288">
          <path
             d="m 2903,1190 h -73 l 58,-12 z m -73,0 58,-12 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11290" />
        </g>
        <g
           id="g11292">
          <path
             d="m 3096,1178 h -66 l 67,-1 z m -66,0 67,-1 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11294" />
        </g>
        <g
           id="g11296">
          <path
             d="m 2888,1178 h -66 l 65,-1 z m -66,0 65,-1 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11298" />
        </g>
        <g
           id="g11300">
          <path
             d="m 3097,1177 h -66 l 72,-15 z m -66,0 72,-15 h -60 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11302" />
        </g>
        <g
           id="g11304">
          <path
             d="m 2887,1177 h -66 l 55,-15 z m -66,0 55,-15 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11306" />
        </g>
        <g
           id="g11308">
          <path
             d="m 3103,1162 h -60 l 63,-8 z m -60,0 63,-8 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11310" />
        </g>
        <g
           id="g11312">
          <path
             d="m 2876,1162 h -61 l 56,-8 z m -61,0 56,-8 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11314" />
        </g>
        <g
           id="g11316">
          <path
             d="m 3106,1154 h -59 l 61,-9 z m -59,0 61,-9 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11318" />
        </g>
        <g
           id="g11320">
          <path
             d="m 2871,1154 h -59 l 54,-9 z m -59,0 54,-9 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11322" />
        </g>
        <g
           id="g11324">
          <path
             d="m 3108,1145 h -56 l 60,-14 z m -56,0 60,-14 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11326" />
        </g>
        <g
           id="g11328">
          <path
             d="m 2866,1145 h -56 l 52,-14 z m -56,0 52,-14 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11330" />
        </g>
        <g
           id="g11332">
          <path
             d="m 3112,1131 h -56 l 56,-5 z m -56,0 56,-5 h -54 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11334" />
        </g>
        <g
           id="g11336">
          <path
             d="m 2862,1131 h -56 l 55,-5 z m -56,0 55,-5 h -55 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11338" />
        </g>
        <g
           id="g11340">
          <path
             d="m 3112,1126 h -54 l 56,-20 z m -54,0 56,-20 h -54 z m 56,-20 h -54 z m -54,0 h 54 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11342" />
        </g>
        <g
           id="g11344">
          <path
             d="m 2861,1126 h -55 l 53,-20 z m -55,0 53,-20 h -54 z m 53,-20 h -54 z m -54,0 h 54 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11346" />
        </g>
        <g
           id="g11348">
          <path
             d="m 3114,1106 h -54 l 52,-19 z m -54,0 52,-19 h -54 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11350" />
        </g>
        <g
           id="g11352">
          <path
             d="m 2859,1106 h -54 l 56,-19 z m -54,0 56,-19 h -55 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11354" />
        </g>
        <g
           id="g11356">
          <path
             d="m 3112,1087 h -54 l 54,-5 z m -54,0 54,-5 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11358" />
        </g>
        <g
           id="g11360">
          <path
             d="m 2861,1087 h -55 l 56,-5 z m -55,0 56,-5 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11362" />
        </g>
        <g
           id="g11364">
          <path
             d="m 3112,1082 h -56 l 52,-14 z m -56,0 52,-14 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11366" />
        </g>
        <g
           id="g11368">
          <path
             d="m 2862,1082 h -56 l 60,-14 z m -56,0 60,-14 h -56 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11370" />
        </g>
        <g
           id="g11372">
          <path
             d="m 3108,1068 h -56 l 54,-9 z m -56,0 54,-9 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11374" />
        </g>
        <g
           id="g11376">
          <path
             d="m 2866,1068 h -56 l 61,-9 z m -56,0 61,-9 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11378" />
        </g>
        <g
           id="g11380">
          <path
             d="m 3106,1059 h -59 l 56,-8 z m -59,0 56,-8 h -60 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11382" />
        </g>
        <g
           id="g11384">
          <path
             d="m 2871,1059 h -59 l 64,-8 z m -59,0 64,-8 h -61 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11386" />
        </g>
        <g
           id="g11388">
          <path
             d="m 3103,1051 h -60 l 54,-15 z m -60,0 54,-15 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11390" />
        </g>
        <g
           id="g11392">
          <path
             d="m 2876,1051 h -61 l 72,-15 z m -61,0 72,-15 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11394" />
        </g>
        <g
           id="g11396">
          <path
             d="m 3097,1036 h -66 l 65,-1 z m -66,0 65,-1 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11398" />
        </g>
        <g
           id="g11400">
          <path
             d="m 2887,1036 h -66 l 67,-1 z m -66,0 67,-1 h -66 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11402" />
        </g>
        <g
           id="g11404">
          <path
             d="m 3096,1035 h -66 l 59,-12 z m -66,0 59,-12 h -74 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11406" />
        </g>
        <g
           id="g11408">
          <path
             d="m 2888,1035 h -66 l 81,-12 z m -66,0 81,-12 h -73 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11410" />
        </g>
        <g
           id="g11412">
          <path
             d="m 3089,1023 h -74 l 69,-7 z m -74,0 69,-7 h -83 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11414" />
        </g>
        <g
           id="g11416">
          <path
             d="m 2903,1023 h -73 l 87,-7 z m -73,0 87,-7 h -83 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11418" />
        </g>
        <g
           id="g11420">
          <path
             d="m 3084,1016 h -83 l 82,-2 z m -83,0 82,-2 h -85 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11422" />
        </g>
        <g
           id="g11424">
          <path
             d="m 2917,1016 h -83 l 87,-2 z m -83,0 87,-2 h -85 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11426" />
        </g>
        <g
           id="g11428">
          <path
             d="m 3083,1014 h -85 l 80,-6 z m -85,0 80,-6 h -99 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11430" />
        </g>
        <g
           id="g11432">
          <path
             d="m 2921,1014 h -85 l 104,-6 z m -85,0 104,-6 h -99 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11434" />
        </g>
        <g
           id="g11436">
          <path
             d="m 3078,1008 h -99 l 97,-2 z m -99,0 97,-2 h -117 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11438" />
        </g>
        <g
           id="g11440">
          <path
             d="m 2940,1008 h -99 l 118,-2 z m -99,0 118,-2 h -117 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11442" />
        </g>
        <g
           id="g11444">
          <path
             d="m 3076,1006 h -117 l 110,-9 z m -117,0 110,-9 h -110 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11446" />
        </g>
        <g
           id="g11448">
          <path
             d="m 2959,1006 h -117 l 117,-9 z m -117,0 117,-9 h -109 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11450" />
        </g>
        <g
           id="g11452">
          <path
             d="m 3069,997 h -110 l 91,-16 z m -110,0 91,-16 h -91 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11454" />
        </g>
        <g
           id="g11456">
          <path
             d="m 2959,997 h -109 l 109,-16 z m -109,0 109,-16 h -91 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11458" />
        </g>
        <g
           id="g11460">
          <path
             d="m 3050,981 h -91 l 70,-12 z m -91,0 70,-12 h -70 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11462" />
        </g>
        <g
           id="g11464">
          <path
             d="m 2959,981 h -91 l 91,-12 z m -91,0 91,-12 h -70 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11466" />
        </g>
        <g
           id="g11468">
          <path
             d="m 3029,969 h -70 l 48,-10 z m -70,0 48,-10 h -48 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11470" />
        </g>
        <g
           id="g11472">
          <path
             d="m 2959,969 h -70 l 70,-10 z m -70,0 70,-10 h -48 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11474" />
        </g>
        <g
           id="g11476">
          <path
             d="m 2935,954 h 24 v -2 z m 24,0 v -2 l 24,2 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11478" />
        </g>
        <g
           id="g11480">
          <path
             d="m 3007,959 h -48 l 24,-5 z m -48,0 24,-5 h -24 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11482" />
        </g>
        <g
           id="g11484">
          <path
             d="m 2959,959 h -48 l 48,-5 z m -48,0 48,-5 h -24 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11486" />
        </g>
        <g
           id="g11488">
          <path
             d="m 2985,1498 33,-6 h -33 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11490" />
        </g>
        <g
           id="g11492">
          <path
             d="m 3018,1492 h -33 l 65,-9 z m -33,0 65,-9 h -65 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11494" />
        </g>
        <g
           id="g11496">
          <path
             d="m 3050,1483 h -65 l 95,-13 z m -65,0 95,-13 h -95 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11498" />
        </g>
        <g
           id="g11500">
          <path
             d="m 3080,1470 h -95 l 124,-16 z m -95,0 124,-16 h -124 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11502" />
        </g>
        <g
           id="g11504">
          <path
             d="m 3109,1454 h -124 l 151,-20 z m -124,0 151,-20 h -151 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11506" />
        </g>
        <g
           id="g11508">
          <path
             d="m 3136,1434 h -151 l 176,-22 z m -151,0 176,-22 h -176 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11510" />
        </g>
        <g
           id="g11512">
          <path
             d="m 3161,1412 h -176 l 197,-26 z m -176,0 197,-26 h -197 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11514" />
        </g>
        <g
           id="g11516">
          <path
             d="m 3182,1386 h -197 l 216,-28 z m -197,0 216,-28 h -216 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11518" />
        </g>
        <g
           id="g11520">
          <path
             d="m 3201,1358 h -216 l 231,-29 z m -216,0 231,-29 h -231 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11522" />
        </g>
        <g
           id="g11524">
          <path
             d="m 3216,1329 h -231 l 243,-32 z m -231,0 243,-32 h -243 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11526" />
        </g>
        <g
           id="g11528">
          <path
             d="m 3228,1297 h -243 l 247,-17 z m -243,0 247,-17 h -247 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11530" />
        </g>
        <g
           id="g11532">
          <path
             d="m 3232,1280 h -247 l 248,-5 z m -247,0 248,-5 h -223 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11534" />
        </g>
        <g
           id="g11536">
          <path
             d="m 3233,1275 h -223 l 225,-10 z m -223,0 225,-10 h -200 z m 225,-10 h -200 z m -200,0 h 200 v 0 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11538" />
        </g>
        <g
           id="g11540">
          <path
             d="m 3235,1265 h -200 l 202,-13 z m -200,0 202,-13 h -179 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11542" />
        </g>
        <g
           id="g11544">
          <path
             d="m 3237,1252 h -179 l 181,-16 z m -179,0 181,-16 h -161 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11546" />
        </g>
        <g
           id="g11548">
          <path
             d="m 3239,1236 h -161 l 161,-4 z m -161,0 161,-4 h -157 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11550" />
        </g>
        <g
           id="g11552">
          <path
             d="m 3239,1232 h -157 l 157,-16 z m -157,0 157,-16 h -143 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11554" />
        </g>
        <g
           id="g11556">
          <path
             d="m 3239,1216 h -143 l 143,-18 z m -143,0 143,-18 h -130 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11558" />
        </g>
        <g
           id="g11560">
          <path
             d="m 3239,1198 h -130 l 130,-3 z m -130,0 130,-3 h -128 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11562" />
        </g>
        <g
           id="g11564">
          <path
             d="m 3239,1195 h -128 l 125,-24 z m -128,0 125,-24 h -113 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11566" />
        </g>
        <g
           id="g11568">
          <path
             d="m 3236,1171 h -113 l 112,-6 z m -113,0 112,-6 h -111 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11570" />
        </g>
        <g
           id="g11572">
          <path
             d="m 3235,1165 h -111 l 107,-19 z m -111,0 107,-19 h -100 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11574" />
        </g>
        <g
           id="g11576">
          <path
             d="m 3231,1146 h -100 l 97,-13 z m -100,0 97,-13 h -96 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11578" />
        </g>
        <g
           id="g11580">
          <path
             d="m 3228,1133 h -96 l 91,-13 z m -96,0 91,-13 h -89 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11582" />
        </g>
        <g
           id="g11584">
          <path
             d="m 3223,1120 h -89 l 82,-18 z m -89,0 82,-18 h -82 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11586" />
        </g>
        <g
           id="g11588">
          <path
             d="m 3216,1102 h -82 l 78,-9 z m -82,0 78,-9 h -78 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11590" />
        </g>
        <g
           id="g11592">
          <path
             d="m 3212,1093 h -78 l 67,-21 z m -78,0 67,-21 h -70 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11594" />
        </g>
        <g
           id="g11596">
          <path
             d="m 3201,1072 h -70 l 67,-5 z m -70,0 67,-5 h -67 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11598" />
        </g>
        <g
           id="g11600">
          <path
             d="m 3198,1067 h -67 l 51,-23 z m -67,0 51,-23 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11602" />
        </g>
        <g
           id="g11604">
          <path
             d="m 3182,1044 h -59 l 58,-2 z m -59,0 58,-2 h -58 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11606" />
        </g>
        <g
           id="g11608">
          <path
             d="m 3181,1042 h -58 l 38,-23 z m -58,0 38,-23 h -50 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11610" />
        </g>
        <g
           id="g11612">
          <path
             d="m 3161,1019 h -50 l 49,-1 z m -50,0 49,-1 h -49 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11614" />
        </g>
        <g
           id="g11616">
          <path
             d="m 3160,1018 h -49 l 26,-21 z m -49,0 26,-21 h -41 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11618" />
        </g>
        <g
           id="g11620">
          <path
             d="m 3137,997 h -41 l 40,-1 z m -41,0 40,-1 h -40 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11622" />
        </g>
        <g
           id="g11624">
          <path
             d="m 3136,996 h -40 l 15,-19 z m -40,0 15,-19 h -33 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11626" />
        </g>
        <g
           id="g11628">
          <path
             d="m 3111,977 h -33 l 31,-1 z m -33,0 31,-1 h -32 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11630" />
        </g>
        <g
           id="g11632">
          <path
             d="m 3109,976 h -32 l 5,-15 z m -32,0 5,-15 h -24 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11634" />
        </g>
        <g
           id="g11636">
          <path
             d="m 3082,961 h -24 l 22,-1 z m -24,0 22,-1 h -24 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11638" />
        </g>
        <g
           id="g11640">
          <path
             d="m 3080,960 h -24 l -5,-12 z m -24,0 -5,-12 h -16 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11642" />
        </g>
        <g
           id="g11644">
          <path
             d="m 3051,948 h -16 l 15,-1 z m -16,0 15,-1 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11646" />
        </g>
        <g
           id="g11648">
          <path
             d="m 3050,947 h -17 l -14,-9 z m -17,0 -14,-9 h -9 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11650" />
        </g>
        <g
           id="g11652">
          <path
             d="m 3010,938 h -1 9 z m -1,0 h 9 l -33,-5 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11654" />
        </g>
        <g
           id="g11656">
          <path
             d="m 3010,938 h 9 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11658" />
        </g>
        <g
           id="g11660">
          <path
             d="m 3285,1261 17,-24 h -17 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11662" />
        </g>
        <g
           id="g11664">
          <path
             d="m 3302,1237 h -17 l 23,-11 z m -17,0 23,-11 h -23 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11666" />
        </g>
        <g
           id="g11668">
          <path
             d="m 3308,1226 h -23 l 31,-16 z m -23,0 31,-16 h -33 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11670" />
        </g>
        <g
           id="g11672">
          <path
             d="m 3316,1210 h -33 l 40,-19 z m -33,0 40,-19 h -42 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11674" />
        </g>
        <g
           id="g11676">
          <path
             d="m 3323,1191 h -42 l 45,-9 z m -42,0 45,-9 h -47 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11678" />
        </g>
        <g
           id="g11680">
          <path
             d="m 3326,1182 h -47 l 53,-25 z m -47,0 53,-25 h -59 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11682" />
        </g>
        <g
           id="g11684">
          <path
             d="m 3332,1157 h -59 l 59,-4 z m -59,0 59,-4 h -60 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11686" />
        </g>
        <g
           id="g11688">
          <path
             d="m 3332,1153 h -60 l 63,-29 z m -60,0 63,-29 h -73 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11690" />
        </g>
        <g
           id="g11692">
          <path
             d="m 3335,1124 h -73 l 73,-1 z m -73,0 73,-1 h -73 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11694" />
        </g>
        <g
           id="g11696">
          <path
             d="m 3335,1123 h -73 l 72,-29 z m -73,0 72,-29 h -85 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11698" />
        </g>
        <g
           id="g11700">
          <path
             d="m 3334,1094 h -85 l 84,-3 z m -85,0 84,-3 h -86 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11702" />
        </g>
        <g
           id="g11704">
          <path
             d="m 3333,1091 h -86 l 82,-26 z m -86,0 82,-26 h -97 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11706" />
        </g>
        <g
           id="g11708">
          <path
             d="m 3329,1065 h -97 l 96,-4 z m -97,0 96,-4 h -98 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11710" />
        </g>
        <g
           id="g11712">
          <path
             d="m 3328,1061 h -98 l 90,-25 z m -98,0 90,-25 h -108 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11714" />
        </g>
        <g
           id="g11716">
          <path
             d="m 3320,1036 h -108 l 107,-4 z m -108,0 107,-4 h -110 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11718" />
        </g>
        <g
           id="g11720">
          <path
             d="m 3319,1032 h -110 l 99,-23 z m -110,0 99,-23 h -120 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11722" />
        </g>
        <g
           id="g11724">
          <path
             d="m 3308,1009 h -120 l 118,-3 z m -120,0 118,-3 h -120 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11726" />
        </g>
        <g
           id="g11728">
          <path
             d="m 3306,1006 h -120 l 107,-22 z m -120,0 107,-22 h -132 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11730" />
        </g>
        <g
           id="g11732">
          <path
             d="m 3293,984 h -132 l 131,-2 z m -132,0 131,-2 h -132 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11734" />
        </g>
        <g
           id="g11736">
          <path
             d="m 3292,982 h -132 l 115,-20 z m -132,0 115,-20 h -144 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11738" />
        </g>
        <g
           id="g11740">
          <path
             d="m 3275,962 h -144 l 143,-1 z m -144,0 143,-1 h -144 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11742" />
        </g>
        <g
           id="g11744">
          <path
             d="m 3274,961 h -144 l 126,-17 z m -144,0 126,-17 h -155 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11746" />
        </g>
        <g
           id="g11748">
          <path
             d="m 3256,944 h -155 l 152,-4 z m -155,0 152,-4 h -159 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11750" />
        </g>
        <g
           id="g11752">
          <path
             d="m 3253,940 h -159 l 143,-11 z m -159,0 143,-11 h -168 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11754" />
        </g>
        <g
           id="g11756">
          <path
             d="m 3237,929 h -168 l 160,-6 z m -168,0 160,-6 h -178 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11758" />
        </g>
        <g
           id="g11760">
          <path
             d="m 3229,923 h -178 l 168,-6 z m -178,0 168,-6 h -183 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11762" />
        </g>
        <g
           id="g11764">
          <path
             d="m 3219,917 h -183 l 169,-8 z m -183,0 169,-8 h -203 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11766" />
        </g>
        <g
           id="g11768">
          <path
             d="m 3205,909 h -203 l 201,-1 z m -203,0 201,-1 h -198 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11770" />
        </g>
        <g
           id="g11772">
          <path
             d="m 3203,908 h -198 l 172,-10 z m -198,0 172,-10 h -148 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11774" />
        </g>
        <g
           id="g11776">
          <path
             d="m 3177,898 h -148 l 146,-1 z m -148,0 146,-1 h -143 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11778" />
        </g>
        <g
           id="g11780">
          <path
             d="m 3175,897 h -143 l 116,-7 z m -143,0 116,-7 h -90 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11782" />
        </g>
        <g
           id="g11784">
          <path
             d="m 3148,890 h -90 89 z m -90,0 h 89 -85 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11786" />
        </g>
        <g
           id="g11788">
          <path
             d="m 3062,890 25,-4 h 31 z m 25,-4 h 31 -1 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11790" />
        </g>
        <g
           id="g11792">
          <path
             d="m 3062,890 h 85 l -29,-4 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path11794" />
        </g>
        <path
           d="m 3647,1370 21,120 h 40 l 17,-6 9,-12 4,-11 2,-17 -5,-29 -8,-17 -8,-11 -14,-12 -18,-5 h -40"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11796" />
        <path
           d="m 3767,1370 21,120 h 75"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11798" />
        <path
           d="m 3778,1432 h 46"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11800" />
        <path
           d="m 3767,1370 h 75"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11802" />
        <path
           d="m 3897,1490 25,-120 66,120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11804" />
        <path
           d="m 3990,1370 21,120 h 75"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11806" />
        <path
           d="m 4001,1432 h 46"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11808" />
        <path
           d="m 3990,1370 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11810" />
        <path
           d="m 4120,1490 -21,-120 h 68"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11812" />
        <path
           d="m 4251,1490 -12,-6 -14,-12 -7,-11 -9,-17 -5,-29 3,-17 3,-11 10,-12 10,-5 h 23 l 12,5 14,12 8,11 8,17 5,29 -2,17 -4,11 -9,12 -11,6 h -23"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11814" />
        <path
           d="m 4322,1370 21,120 h 51 l 16,-6 5,-6 4,-11 -3,-17 -8,-12 -7,-6 -18,-5 h -51"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11816" />
        <path
           d="m 4442,1370 21,120 24,-120 67,120 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11818" />
        <path
           d="m 4579,1370 21,120 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11820" />
        <path
           d="m 4590,1432 h 45"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11822" />
        <path
           d="m 4579,1370 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11824" />
        <path
           d="m 4687,1370 21,120 59,-120 21,120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11826" />
        <path
           d="m 4874,1490 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11828" />
        <path
           d="m 4834,1490 h 80"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11830" />
        <path
           d="m 5122,1472 -9,12 -16,6 h -23 l -18,-6 -14,-12 -2,-11 4,-11 5,-6 10,-6 33,-11 10,-6 5,-6 3,-11 -3,-17 -13,-12 -18,-5 h -23 l -16,5 -10,12"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11832" />
        <path
           d="m 5139,1370 21,120 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11834" />
        <path
           d="m 5150,1432 h 45"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11836" />
        <path
           d="m 5139,1370 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11838" />
        <path
           d="m 5247,1370 21,120 h 52 l 16,-6 5,-6 3,-11 -2,-12 -7,-11 -7,-6 -18,-6 h -52"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11840" />
        <path
           d="m 5298,1432 29,-62"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11842" />
        <path
           d="m 5388,1490 25,-120 67,120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11844" />
        <path
           d="m 5481,1370 22,120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11846" />
        <path
           d="m 5629,1461 -4,11 -9,12 -11,6 h -22 l -13,-6 -13,-12 -8,-11 -9,-17 -5,-29 3,-17 4,-11 9,-12 10,-5 h 23 l 13,5 13,12 8,11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11848" />
        <path
           d="m 5647,1370 21,120 h 75"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11850" />
        <path
           d="m 5658,1432 h 46"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11852" />
        <path
           d="m 5647,1370 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11854" />
        <path
           d="m 5854,1472 -10,12 -16,6 h -23 l -18,-6 -13,-12 -2,-11 4,-11 4,-6 11,-6 32,-11 10,-6 5,-6 4,-11 -3,-17 -14,-12 -18,-5 h -23 l -16,5 -9,12"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11856" />
        <path
           d="m 5979,1370 21,120 h 40 l 16,-6 9,-12 4,-11 3,-17 -5,-29 -9,-17 -8,-11 -13,-12 -18,-5 h -40"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11858" />
        <path
           d="m 6099,1370 21,120 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11860" />
        <path
           d="m 6110,1432 h 45"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11862" />
        <path
           d="m 6099,1370 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11864" />
        <path
           d="m 6207,1370 21,120 h 52 l 16,-6 5,-6 3,-11 -3,-17 -7,-12 -7,-6 -18,-5 h -52"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11866" />
        <path
           d="m 6327,1370 67,120 25,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11868" />
        <path
           d="m 6351,1410 h 57"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11870" />
        <path
           d="m 6453,1370 21,120 h 51 l 17,-6 4,-6 4,-11 -2,-12 -8,-11 -6,-6 -19,-6 h -51"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11872" />
        <path
           d="m 6504,1432 29,-62"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11874" />
        <path
           d="m 6634,1490 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11876" />
        <path
           d="m 6594,1490 h 80"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11878" />
        <path
           d="m 6676,1370 21,120 24,-120 67,120 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11880" />
        <path
           d="m 6813,1370 21,120 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11882" />
        <path
           d="m 6824,1432 h 46"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11884" />
        <path
           d="m 6813,1370 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11886" />
        <path
           d="m 6921,1370 22,120 58,-120 22,120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11888" />
        <path
           d="m 7108,1490 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11890" />
        <path
           d="m 7068,1490 h 80"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11892" />
        <path
           d="m 3745,1118 -9,11 -16,6 h -23 l -18,-6 -14,-11 -2,-11 4,-12 5,-6 10,-5 32,-12 11,-5 5,-6 3,-12 -3,-17 -13,-11 -18,-6 h -23 l -16,6 -10,11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11894" />
        <path
           d="m 3762,1015 66,120 25,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11896" />
        <path
           d="m 3786,1055 h 57"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11898" />
        <path
           d="m 3887,1015 21,120 59,-120 21,120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11900" />
        <path
           d="m 4122,1015 21,120 h 40 l 16,-6 9,-11 4,-11 3,-18 -5,-28 -9,-17 -8,-12 -13,-11 -18,-6 h -40"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11902" />
        <path
           d="m 4242,1015 21,120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11904" />
        <path
           d="m 4287,1015 21,120 h 75"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11906" />
        <path
           d="m 4298,1078 h 46"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11908" />
        <path
           d="m 4287,1015 h 75"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11910" />
        <path
           d="m 4498,1107 -4,11 -9,11 -11,6 h -23 l -12,-6 -14,-11 -7,-11 -9,-18 -5,-28 3,-17 3,-12 10,-11 10,-6 h 23 l 12,6 14,11 8,12 3,17 h -29"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11912" />
        <path
           d="m 4571,1135 -12,-6 -14,-11 -7,-11 -9,-18 -5,-28 3,-17 3,-12 10,-11 10,-6 h 23 l 12,6 14,11 8,12 8,17 5,28 -2,18 -4,11 -9,11 -11,6 h -23"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11914" />
        <path
           d="m 4654,1021 -7,-6 -4,6 6,6 5,-6 -2,-12 -8,-11 -7,-6"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11916" />
        <path
           d="m 4909,1107 -4,11 -9,11 -10,6 h -23 l -13,-6 -13,-11 -8,-11 -9,-18 -5,-28 3,-17 4,-12 9,-11 10,-6 h 23 l 13,6 13,11 8,12"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11918" />
        <path
           d="m 4927,1015 67,120 25,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11920" />
        <path
           d="m 4951,1055 h 58"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11922" />
        <path
           d="m 5250,1095 -9,-17 -13,-11 -18,-6 h -6 l -16,6 -10,11 -2,17 1,6 8,17 14,11 18,6 h 6 l 16,-6 9,-11 2,-23 -5,-28 -11,-29 -14,-17 -19,-6 h -11 l -16,6 -4,11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11924" />
        <path
           d="m 5298,1107 1,5 7,12 7,5 12,6 h 23 l 11,-6 4,-5 4,-12 -2,-11 -8,-12 -14,-17 -67,-57 h 80"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11926" />
        <path
           d="m 5407,1112 13,6 20,17 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11928" />
        <path
           d="m 5537,1135 -18,-6 -15,-17 -10,-28 -3,-17 v -29 l 9,-17 16,-6 h 11 l 18,6 15,17 11,29 3,17 -1,28 -9,17 -16,6 h -11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11930" />
        <path
           d="m 5613,1112 12,6 20,17 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11932" />
        <path
           d="m 5696,1067 h 103"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11934" />
        <path
           d="m 5893,1015 21,120 -71,-80 h 85"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11936" />
        <path
           d="m 5967,1112 13,6 20,17 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11938" />
        <path
           d="m 6131,1135 h -57 l -15,-51 7,5 18,6 h 17 l 16,-6 10,-11 2,-17 -2,-12 -8,-17 -14,-11 -18,-6 h -17 l -16,6 -5,6 -4,11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11940" />
        <path
           d="m 6245,1135 h -57 l -14,-51 6,5 18,6 h 18 l 16,-6 9,-11 3,-17 -2,-12 -9,-17 -13,-11 -19,-6 h -17 l -16,6 -5,6 -3,11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11942" />
        <path
           d="m 3664,1290 13,5 20,17 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11944" />
        <path
           d="m 3761,1284 1,6 7,11 7,6 12,5 h 23 l 11,-5 4,-6 4,-11 -2,-12 -8,-11 -14,-17 -67,-58 h 80"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11946" />
        <path
           d="m 3875,1284 1,6 8,11 6,6 13,5 h 23 l 10,-5 5,-6 3,-11 -2,-12 -7,-11 -15,-17 -67,-58 h 80"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11948" />
        <path
           d="m 3989,1284 1,6 8,11 7,6 12,5 h 23 l 10,-5 5,-6 4,-11 -2,-12 -8,-11 -15,-17 -67,-58 h 80"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11950" />
        <path
           d="m 4207,1290 13,5 20,17 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11952" />
        <path
           d="m 4380,1295 -10,12 -16,5 h -23 l -18,-5 -13,-12 -2,-11 3,-12 5,-5 10,-6 33,-11 10,-6 5,-6 4,-11 -3,-17 -14,-12 -18,-6 h -23 l -16,6 -9,12"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11954" />
        <path
           d="m 4457,1312 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11956" />
        <path
           d="m 4417,1312 h 80"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11958" />
        <path
           d="m 4607,1192 67,120 25,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11960" />
        <path
           d="m 4631,1232 h 58"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11962" />
        <path
           d="m 4754,1312 25,-120 67,120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11964" />
        <path
           d="m 4847,1192 21,120 h 75"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11966" />
        <path
           d="m 4858,1255 h 46"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11968" />
        <path
           d="m 4847,1192 h 74"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11970" />
        <path
           d="m 3734,941 -4,11 -16,6 h -11 l -18,-6 -15,-17 -11,-28 -5,-29 2,-23 9,-11 17,-6 h 5 l 18,6 14,11 9,17 1,6 -3,17 -10,12 -16,5 h -5 l -19,-5 -13,-12 -9,-17"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11972" />
        <path
           d="m 3779,935 12,6 20,17 -21,-120"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11974" />
        <path
           d="m 3941,918 -8,-17 -14,-12 -18,-5 h -6 l -16,5 -9,12 -3,17 1,6 9,17 13,11 18,6 h 6 l 16,-6 10,-11 1,-23 -5,-29 -10,-28 -15,-17 -18,-6 h -11 l -17,6 -3,11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11976" />
        <path
           d="m 3976,889 h 103"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11978" />
        <path
           d="m 4173,838 21,120 -71,-80 h 86"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11980" />
        <path
           d="m 4287,838 21,120 -71,-80 h 86"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11982" />
        <path
           d="m 4431,941 -4,11 -16,6 h -11 l -18,-6 -15,-17 -11,-28 -5,-29 2,-23 10,-11 16,-6 h 5 l 19,6 13,11 9,17 1,6 -3,17 -9,12 -17,5 h -5 l -18,-5 -14,-12 -9,-17"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11984" />
        <path
           d="m 4468,889 h 103"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11986" />
        <path
           d="m 4697,958 h -57 l -15,-51 7,5 18,6 h 17 l 16,-6 10,-11 2,-17 -2,-12 -8,-17 -14,-11 -18,-6 h -17 l -16,6 -5,5 -4,12"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11988" />
        <path
           d="m 4777,958 -18,-6 -15,-17 -10,-28 -3,-18 v -28 l 9,-17 16,-6 h 11 l 18,6 15,17 11,28 3,18 -1,28 -9,17 -16,6 h -11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11990" />
        <path
           d="m 4891,958 -18,-6 -14,-17 -11,-28 -3,-18 1,-28 8,-17 16,-6 h 11 l 19,6 14,17 11,28 3,18 -1,28 -8,17 -16,6 h -12"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11992" />
        <path
           d="m 5005,958 -18,-6 -14,-17 -11,-28 -3,-18 1,-28 8,-17 16,-6 h 12 l 18,6 14,17 11,28 3,18 -1,28 -8,17 -16,6 h -12"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11994" />
        <path
           d="m 4278,211 -3,12 -10,11 -10,6 h -23 l -12,-6 -13,-11 -8,-12 -8,-16 -5,-29 2,-16 4,-12 9,-11 11,-6 h 22 l 12,6 14,11 7,12"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11996" />
        <path
           d="m 4351,240 -13,-6 -13,-11 -7,-12 -9,-16 -5,-29 3,-16 3,-12 10,-11 10,-6 h 22 l 13,6 13,11 7,12 9,16 5,29 -3,16 -3,12 -10,11 -10,6 h -22"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path11998" />
        <path
           d="m 4420,121 21,119 58,-119 20,119"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12000" />
        <path
           d="m 4640,223 -9,11 -16,6 h -22 l -18,-6 -14,-11 -2,-12 4,-11 5,-5 10,-6 32,-11 10,-6 5,-6 3,-11 -3,-17 -13,-11 -18,-6 h -22 l -16,6 -9,11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12002" />
        <path
           d="M 4716,240 4695,121"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12004" />
        <path
           d="m 4677,240 h 79"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12006" />
        <path
           d="m 4757,121 21,119 h 51 l 16,-6 4,-6 4,-11 -2,-11 -8,-11 -6,-6 -18,-6 h -51"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12008" />
        <path
           d="m 4808,183 28,-62"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12010" />
        <path
           d="m 4896,240 -15,-85 3,-17 9,-11 16,-6 h 11 l 18,6 14,11 8,17 15,85"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12012" />
        <path
           d="m 5099,211 -3,12 -9,11 -11,6 h -22 l -12,-6 -14,-11 -7,-12 -9,-16 -5,-29 3,-16 3,-12 10,-11 10,-6 h 22 l 13,6 13,11 8,12"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12014" />
        <path
           d="M 5178,240 5157,121"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12016" />
        <path
           d="m 5138,240 h 79"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12018" />
        <path
           d="m 5219,121 20,119"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12020" />
        <path
           d="m 5318,240 -12,-6 -13,-11 -8,-12 -9,-16 -4,-29 2,-16 4,-12 9,-11 10,-6 h 23 l 12,6 13,11 8,12 9,16 5,29 -3,16 -4,12 -9,11 -10,6 h -23"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12022" />
        <path
           d="m 5387,121 21,119 58,-119 21,119"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12024" />
        <path
           d="m 5618,121 21,119 h 50 l 16,-6 5,-6 4,-11 -3,-17 -8,-11 -7,-6 -17,-5 h -51"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12026" />
        <path
           d="m 5757,240 -21,-119 h 68"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12028" />
        <path
           d="m 5832,121 66,119 24,-119"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12030" />
        <path
           d="m 5856,161 h 56"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12032" />
        <path
           d="m 5956,121 20,119 58,-119 21,119"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12034" />
        <path
           d="m 6186,121 21,119 h 39 l 16,-6 10,-11 3,-12 3,-16 -5,-29 -9,-16 -7,-12 -14,-11 -17,-6 h -40"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12036" />
        <path
           d="m 6401,223 -9,11 -16,6 h -23 l -18,-6 -13,-11 -2,-12 4,-11 4,-5 11,-6 31,-11 11,-6 4,-6 4,-11 -3,-17 -13,-11 -18,-6 h -23 l -15,6 -10,11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12038" />
        <path
           d="m 6426,172 h 101"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12040" />
        <path
           d="m 6595,240 h 62 l -42,-45 h 17 l 10,-6 5,-6 3,-17 -2,-11 -9,-17 -13,-11 -18,-6 h -17 l -16,6 -4,6 -4,11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12042" />
        <path
           d="m 6692,217 13,6 20,17 -21,-119"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12044" />
        <path
           d="m 6786,240 h 79 l -77,-119"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12046" />
        <path
           d="m 6965,200 -8,-17 -14,-11 -18,-6 h -5 l -16,6 -9,11 -3,17 1,6 9,17 13,11 18,6 h 5 l 16,-6 9,-11 2,-23 -5,-28 -10,-28 -15,-17 -18,-6 h -11 l -16,6 -3,11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12048" />
        <path
           d="m 7269,262 -14,-11 -14,-17 -15,-23 -11,-28 -4,-22 1,-28 7,-23 9,-17 9,-11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12050" />
        <path
           d="m 7300,217 12,6 20,17 -21,-119"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12052" />
        <path
           d="m 7395,211 1,6 7,11 7,6 12,6 h 23 l 10,-6 4,-6 4,-11 -2,-11 -7,-11 -15,-17 -66,-57 h 79"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12054" />
        <path
           d="M 7612,262 7479,82"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12056" />
        <path
           d="m 7695,223 -4,11 -16,6 h -11 l -18,-6 -14,-17 -11,-28 -5,-28 2,-23 9,-11 16,-6 h 6 l 18,6 13,11 8,17 1,6 -2,17 -9,11 -16,6 h -6 l -18,-6 -13,-11 -9,-17"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12058" />
        <path
           d="M 7848,262 7715,82"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12060" />
        <path
           d="m 7867,211 1,6 8,11 6,6 13,6 h 22 l 10,-6 5,-6 4,-11 -2,-11 -8,-11 -14,-17 -66,-57 h 78"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12062" />
        <path
           d="m 8013,240 -18,-6 -14,-17 -11,-28 -3,-17 1,-28 8,-17 16,-6 h 11 l 18,6 14,17 11,28 3,17 -1,28 -8,17 -16,6 h -11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12064" />
        <path
           d="m 8092,211 1,6 8,11 6,6 13,6 h 22 l 10,-6 5,-6 4,-11 -2,-11 -8,-11 -14,-17 -66,-57 h 78"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12066" />
        <path
           d="m 8200,217 12,6 20,17 -21,-119"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12068" />
        <path
           d="m 8298,262 9,-11 9,-17 7,-23 v -28 l -3,-22 -11,-28 -15,-23 -15,-17 -13,-11"
           style="fill:none;stroke:#0000ff;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12070" />
        <g
           id="g12072">
          <path
             d="m 10953,1786 h -12 l 12,-1321 z m -12,0 12,-1321 h -12 z"
             style="fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:#0000ff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12074" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.83670722,0,-0.17361286,-0.98481398,7629,1168)"
           style="font-variant:normal;font-weight:normal;font-size:168.895px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12078"><tspan
             x="0 95.71093 199.31406 271.06137 310.95288 414.55603 526.19489 566.08636"
             y="0"
             sodipodi:role="line"
             id="tspan12076">PRJ NO: </tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(0.83670722,0,-0.17361286,-0.98481398,8226,1168)"
           style="font-variant:normal;font-weight:normal;font-size:168.895px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12082"><tspan
             x="0 79.78302 159.56604 239.34906 319.13208 398.9151 478.69812"
             y="0"
             sodipodi:role="line"
             id="tspan12080">1067219</tspan></text>
        <g
           id="g12084">
          <path
             d="m 12185,1780 v 11 l -5742,-11 z m 0,11 -5742,-11 v 11 z"
             style="fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:#0000ff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12086" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.83670722,0,-0.17361286,-0.98481398,7596,591)"
           style="font-variant:normal;font-weight:normal;font-size:168.895px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12090"><tspan
             x="0 95.71093 199.31406 295.02499 390.7359 478.41113"
             y="0"
             sodipodi:role="line"
             id="tspan12088">SHEET </tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(0.83670722,0,-0.17361286,-0.98481398,8107,591)"
           style="font-variant:normal;font-weight:normal;font-size:168.895px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12094"><tspan
             x="0"
             y="0"
             id="tspan12092">6</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(0.83670722,0,-0.17361286,-0.98481398,8224.2857,591)"
           style="font-variant:normal;font-weight:normal;font-size:168.895px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12098"><tspan
             x="0 111.63883 199.31406"
             y="0"
             sodipodi:role="line"
             id="tspan12096">OF </tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(0.83670722,0,-0.17361286,-0.98481398,8460,591)"
           style="font-variant:normal;font-weight:normal;font-size:168.895px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12102"><tspan
             x="0"
             y="0"
             id="tspan12100">6</tspan></text>
        <g
           id="g12104">
          <path
             d="m 12185,1780 v 11 L 445,1780 Z m 0,11 -11740,-11 v 11 z"
             style="fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:#0000ff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12106" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.83670722,0,-0.17361286,-0.98481398,7611,880)"
           style="font-variant:normal;font-weight:normal;font-size:168.895px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12110"><tspan
             x="0 95.71093 215.24196 302.91721 342.80872 446.41183 558.05066 597.9422"
             y="0"
             sodipodi:role="line"
             id="tspan12108">PMT NO: </tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(0.83670722,0,-0.17361286,-0.98481398,8240,880)"
           style="font-variant:normal;font-weight:normal;font-size:168.895px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12114"><tspan
             x="0 79.78302 159.56604 239.34906 319.13208 398.9151 478.69812"
             y="0"
             sodipodi:role="line"
             id="tspan12112">3171537</tspan></text>
        <g
           id="g12116">
          <path
             d="m 8640,3710 h -12 l 12,-1924 z m -12,0 12,-1924 h -12 z"
             style="fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:#0000ff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12118" />
        </g>
        <g
           id="g12120">
          <path
             d="m 7337,1787 h -12 l 12,-1320 z m -12,0 12,-1320 h -12 z"
             style="fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:#0000ff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12122" />
        </g>
        <g
           id="g12124">
          <path
             d="m 12204,3704 v 12 l -3570,-12 z m 0,12 -3570,-12 v 12 z"
             style="fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:#0000ff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12126" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.78765885,0,-0.17361286,-0.98481398,11297,985)"
           style="font-variant:normal;font-weight:normal;font-size:394.104px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12130"><tspan
             x="0 227.57883 402.83344"
             y="0"
             sodipodi:role="line"
             id="tspan12128">C02</tspan></text>
        <path
           d="m 1626,3847 v -86 l 5,-17 12,-11 17,-6 h 11 l 18,6 11,11 6,17 v 86"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12132" />
        <path
           d="M 1791,3847 V 3727"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12134" />
        <path
           d="m 1751,3847 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12136" />
        <path
           d="m 1854,3727 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12138" />
        <path
           d="m 1900,3847 v -120 h 69"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12140" />
        <path
           d="m 1997,3727 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12142" />
        <path
           d="M 2083,3847 V 3727"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12144" />
        <path
           d="m 2043,3847 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12146" />
        <path
           d="m 2146,3847 45,-57 46,57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12148" />
        <path
           d="m 2191,3790 v -63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12150" />
        <path
           d="m 2454,3818 -6,12 -11,11 -11,6 h -23 l -12,-6 -11,-11 -6,-12 -5,-17 v -28 l 5,-17 6,-12 11,-11 12,-6 h 23 l 11,6 11,11 6,12"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12152" />
        <path
           d="m 2488,3727 v 120 h 52 l 17,-6 6,-5 5,-12 v -11 l -5,-12 -6,-5 -17,-6 h -52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12154" />
        <path
           d="m 2528,3790 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12156" />
        <path
           d="m 2643,3847 -12,-6 -11,-11 -6,-12 -6,-17 v -28 l 6,-17 6,-12 11,-11 12,-6 h 23 l 11,6 11,11 6,12 6,17 v 28 l -6,17 -6,12 -11,11 -11,6 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12158" />
        <path
           d="m 2814,3830 -11,11 -17,6 h -23 l -17,-6 -12,-11 v -12 l 6,-11 6,-6 11,-5 34,-12 12,-6 5,-5 6,-12 v -17 l -11,-11 -17,-6 h -23 l -17,6 -12,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12160" />
        <path
           d="m 2928,3830 -11,11 -17,6 h -23 l -17,-6 -12,-11 v -12 l 6,-11 6,-6 11,-5 35,-12 11,-6 6,-5 5,-12 v -17 l -11,-11 -17,-6 h -23 l -17,6 -12,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12162" />
        <path
           d="m 2963,3727 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12164" />
        <path
           d="m 3008,3727 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12166" />
        <path
           d="m 3220,3818 -6,12 -11,11 -12,6 h -23 l -11,-6 -11,-11 -6,-12 -6,-17 v -28 l 6,-17 6,-12 11,-11 11,-6 h 23 l 12,6 11,11 6,12 v 17 h -29"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12168" />
        <path
           d="m 3363,3727 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12170" />
        <path
           d="m 3408,3727 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12172" />
        <path
           d="m 3534,3727 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12174" />
        <path
           d="m 3534,3790 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12176" />
        <path
           d="m 3671,3847 -11,-6 -12,-11 -5,-12 -6,-17 v -28 l 6,-17 5,-12 12,-11 11,-6 h 23 l 12,6 11,11 6,12 5,17 v 28 l -5,17 -6,12 -11,11 -12,6 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12178" />
        <path
           d="m 3763,3727 v 120 h 51 l 17,-6 6,-5 6,-12 v -11 l -6,-12 -6,-5 -17,-6 h -51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12180" />
        <path
           d="m 3803,3790 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12182" />
        <path
           d="m 3883,3727 v 120 l 45,-120 46,120 v -120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12184" />
        <path
           d="m 4020,3727 46,120 45,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12186" />
        <path
           d="m 4037,3767 h 57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12188" />
        <path
           d="M 4186,3847 V 3727"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12190" />
        <path
           d="m 4146,3847 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12192" />
        <path
           d="m 4248,3727 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12194" />
        <path
           d="m 4328,3847 -11,-6 -11,-11 -6,-12 -6,-17 v -28 l 6,-17 6,-12 11,-11 11,-6 h 23 l 12,6 11,11 6,12 6,17 v 28 l -6,17 -6,12 -11,11 -12,6 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12196" />
        <path
           d="m 4420,3727 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12198" />
        <path
           d="m 915,3483 v -86 l 6,-17 11,-11 17,-6 h 12 l 17,6 11,11 6,17 v 86"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12200" />
        <path
           d="M 1081,3483 V 3363"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12202" />
        <path
           d="m 1041,3483 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12204" />
        <path
           d="m 1144,3363 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12206" />
        <path
           d="m 1189,3483 v -120 h 69"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12208" />
        <path
           d="m 1286,3363 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12210" />
        <path
           d="M 1372,3483 V 3363"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12212" />
        <path
           d="m 1332,3483 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12214" />
        <path
           d="m 1435,3483 46,-57 45,57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12216" />
        <path
           d="m 1481,3426 v -63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12218" />
        <path
           d="m 824,3254 -6,12 -12,11 -11,6 h -23 l -11,-6 -12,-11 -5,-12 -6,-17 v -28 l 6,-17 5,-12 12,-11 11,-6 h 23 l 11,6 12,11 6,12"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12220" />
        <path
           d="m 858,3163 v 120 h 51 l 17,-6 6,-5 6,-12 v -11 l -6,-12 -6,-5 -17,-6 h -51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12222" />
        <path
           d="m 898,3226 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12224" />
        <path
           d="m 1012,3283 -11,-6 -12,-11 -5,-12 -6,-17 v -28 l 6,-17 5,-12 12,-11 11,-6 h 23 l 11,6 12,11 6,12 5,17 v 28 l -5,17 -6,12 -12,11 -11,6 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12226" />
        <path
           d="m 1184,3266 -12,11 -17,6 h -23 l -17,-6 -11,-11 v -12 l 5,-11 6,-6 11,-5 35,-12 11,-6 6,-5 6,-12 v -17 l -12,-11 -17,-6 h -23 l -17,6 -11,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12228" />
        <path
           d="m 1298,3266 -12,11 -17,6 h -23 l -17,-6 -11,-11 v -12 l 6,-11 5,-6 12,-5 34,-12 11,-6 6,-5 6,-12 v -17 l -12,-11 -17,-6 h -23 l -17,6 -11,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12230" />
        <path
           d="m 1332,3163 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12232" />
        <path
           d="m 1378,3163 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12234" />
        <path
           d="m 1589,3254 -5,12 -12,11 -11,6 h -23 l -12,-6 -11,-11 -6,-12 -5,-17 v -28 l 5,-17 6,-12 11,-11 12,-6 h 23 l 11,6 12,11 5,12 v 17 h -28"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12236" />
        <path
           d="m 1704,3266 -12,11 -17,6 h -23 l -17,-6 -11,-11 v -12 l 5,-11 6,-6 11,-5 35,-12 11,-6 6,-5 6,-12 v -17 l -12,-11 -17,-6 h -23 l -17,6 -11,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12238" />
        <path
           d="m 2519,3383 v -86 l 6,-17 11,-11 17,-6 h 12 l 17,6 11,11 6,17 v 86"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12240" />
        <path
           d="M 2685,3383 V 3263"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12242" />
        <path
           d="m 2645,3383 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12244" />
        <path
           d="m 2748,3263 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12246" />
        <path
           d="m 2793,3383 v -120 h 69"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12248" />
        <path
           d="m 2890,3263 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12250" />
        <path
           d="M 2976,3383 V 3263"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12252" />
        <path
           d="m 2936,3383 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12254" />
        <path
           d="m 3039,3383 46,-57 45,57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12256" />
        <path
           d="m 3085,3326 v -63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12258" />
        <path
           d="m 3348,3354 -6,12 -12,11 -11,6 h -23 l -11,-6 -12,-11 -5,-12 -6,-17 v -28 l 6,-17 5,-12 12,-11 11,-6 h 23 l 11,6 12,11 6,12"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12260" />
        <path
           d="m 3382,3263 v 120 h 51 l 17,-6 6,-5 6,-12 v -11 l -6,-12 -6,-5 -17,-6 h -51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12262" />
        <path
           d="m 3422,3326 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12264" />
        <path
           d="m 3536,3383 -11,-6 -12,-11 -5,-12 -6,-17 v -28 l 6,-17 5,-12 12,-11 11,-6 h 23 l 11,6 12,11 6,12 5,17 v 28 l -5,17 -6,12 -12,11 -11,6 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12266" />
        <path
           d="m 3708,3366 -12,11 -17,6 h -23 l -17,-6 -11,-11 v -12 l 5,-11 6,-6 11,-5 35,-12 11,-6 6,-5 6,-12 v -17 l -12,-11 -17,-6 h -23 l -17,6 -11,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12268" />
        <path
           d="m 3822,3366 -12,11 -17,6 h -23 l -17,-6 -11,-11 v -12 l 6,-11 5,-6 12,-5 34,-12 11,-6 6,-5 6,-12 v -17 l -12,-11 -17,-6 h -23 l -17,6 -11,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12270" />
        <path
           d="m 3856,3263 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12272" />
        <path
           d="m 3902,3263 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12274" />
        <path
           d="m 4113,3354 -5,12 -12,11 -11,6 h -23 l -12,-6 -11,-11 -6,-12 -5,-17 v -28 l 5,-17 6,-12 11,-11 12,-6 h 23 l 11,6 12,11 5,12 v 17 h -28"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12276" />
        <path
           d="m 4256,3263 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12278" />
        <path
           d="m 4416,3383 -11,-6 -12,-11 -5,-12 -6,-17 v -28 l 6,-17 5,-12 12,-11 11,-6 h 23 l 11,6 12,11 6,12 5,17 v 28 l -5,17 -6,12 -12,11 -11,6 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12280" />
        <path
           d="M 4548,3383 V 3263"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12282" />
        <path
           d="m 4508,3383 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12284" />
        <path
           d="m 4610,3263 v 120 h 75"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12286" />
        <path
           d="m 4610,3326 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12288" />
        <path
           d="m 4610,3263 h 75"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12290" />
        <path
           d="m 4799,3366 -11,11 -18,6 h -22 l -18,-6 -11,-11 v -12 l 6,-11 5,-6 12,-5 34,-12 12,-6 5,-5 6,-12 v -17 l -11,-11 -18,-6 h -22 l -18,6 -11,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12292" />
        <path
           d="m 1095,2596 29,-120 28,120 29,-120 28,120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12294" />
        <path
           d="m 1238,2556 -6,-6 6,-5 6,5 -6,6"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12296" />
        <path
           d="m 1238,2488 -6,-6 6,-6 6,6 -6,6"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12298" />
        <path
           d="m 1318,2573 11,6 17,17 v -120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12300" />
        <path
           d="m 1889,2876 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12302" />
        <path
           d="m 1889,2939 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12304" />
        <path
           d="m 1889,2876 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12306" />
        <path
           d="m 1998,2876 80,120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12308" />
        <path
           d="m 1998,2996 80,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12310" />
        <path
           d="m 2112,2876 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12312" />
        <path
           d="m 2238,2979 -12,11 -17,6 h -23 l -17,-6 -11,-11 v -11 l 5,-12 6,-6 11,-5 35,-12 11,-5 6,-6 6,-12 v -17 l -12,-11 -17,-6 h -23 l -17,6 -11,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12314" />
        <path
           d="M 2312,2996 V 2876"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12316" />
        <path
           d="m 2272,2996 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12318" />
        <path
           d="m 2375,2876 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12320" />
        <path
           d="m 2420,2876 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12322" />
        <path
           d="m 2632,2968 -6,11 -11,11 -12,6 h -23 l -11,-6 -11,-11 -6,-11 -6,-18 v -28 l 6,-17 6,-12 11,-11 11,-6 h 23 l 12,6 11,11 6,12 v 17 h -29"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12324" />
        <path
           d="m 2775,2973 11,6 17,17 v -120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12326" />
        <path
           d="m 2877,3013 -5,-5 -6,5 6,6 5,-6 v -11 l -5,-12 -6,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12328" />
        <path
           d="m 2912,3013 -6,-5 -6,5 6,6 6,-6 v -11 l -6,-12 -6,-5"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12330" />
        <path
           d="m 3060,2996 29,-120 28,120 29,-120 29,120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12332" />
        <path
           d="m 3197,2876 46,120 46,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12334" />
        <path
           d="m 3215,2916 h 57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12336" />
        <path
           d="M 3363,2996 V 2876"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12338" />
        <path
           d="m 3323,2996 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12340" />
        <path
           d="m 3426,2876 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12342" />
        <path
           d="m 3426,2939 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12344" />
        <path
           d="m 3426,2876 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12346" />
        <path
           d="m 3535,2876 v 120 h 51 l 17,-6 6,-5 6,-12 v -11 l -6,-12 -6,-5 -17,-6 h -51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12348" />
        <path
           d="m 3575,2939 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12350" />
        <path
           d="m 3763,2996 v -120 h 69"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12352" />
        <path
           d="m 3860,2876 46,120 46,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12354" />
        <path
           d="m 3877,2916 h 58"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12356" />
        <path
           d="M 4026,2996 V 2876"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12358" />
        <path
           d="m 3986,2996 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12360" />
        <path
           d="m 4089,2876 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12362" />
        <path
           d="m 4089,2939 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12364" />
        <path
           d="m 4089,2876 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12366" />
        <path
           d="m 4197,2876 v 120 h 52 l 17,-6 6,-5 5,-12 v -11 l -5,-12 -6,-5 -17,-6 h -52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12368" />
        <path
           d="m 4237,2939 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12370" />
        <path
           d="m 4317,2876 46,120 46,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12372" />
        <path
           d="m 4335,2916 h 57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12374" />
        <path
           d="m 4443,2996 v -120 h 69"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12376" />
        <path
           d="m 4649,2876 v 120 h 51 l 17,-6 6,-5 6,-12 v -17 l -6,-11 -6,-6 -17,-6 h -51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12378" />
        <path
           d="m 4769,2876 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12380" />
        <path
           d="m 4769,2939 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12382" />
        <path
           d="m 4769,2876 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12384" />
        <path
           d="m 4877,2876 v 120 h 52 l 17,-6 6,-5 5,-12 v -11 l -5,-12 -6,-5 -17,-6 h -52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12386" />
        <path
           d="m 4917,2939 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12388" />
        <path
           d="m 1889,2676 v 120 h 40 l 17,-6 12,-11 5,-11 6,-18 v -28 l -6,-17 -5,-12 -12,-11 -17,-6 h -40"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12390" />
        <path
           d="m 2009,2676 v 120 h 51 l 18,-6 5,-5 6,-12 v -11 l -6,-12 -5,-5 -18,-6 h -51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12392" />
        <path
           d="m 2049,2739 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12394" />
        <path
           d="m 2129,2676 46,120 45,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12396" />
        <path
           d="m 2146,2716 h 57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12398" />
        <path
           d="m 2255,2796 28,-120 29,120 28,-120 29,120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12400" />
        <path
           d="m 2392,2676 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12402" />
        <path
           d="m 2438,2676 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12404" />
        <path
           d="m 2649,2768 -6,11 -11,11 -12,6 h -22 l -12,-6 -11,-11 -6,-11 -6,-18 v -28 l 6,-17 6,-12 11,-11 12,-6 h 22 l 12,6 11,11 6,12 v 17 h -29"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12406" />
        <path
           d="m 2792,2676 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12408" />
        <path
           d="m 2952,2796 -12,-6 -11,-11 -6,-11 -6,-18 v -28 l 6,-17 6,-12 11,-11 12,-6 h 23 l 11,6 11,11 6,12 6,17 v 28 l -6,18 -6,11 -11,11 -11,6 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12410" />
        <path
           d="m 3049,2688 -6,-6 6,-6 6,6"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12412" />
        <path
           d="m 3220,2796 h 63 l -34,-46 h 17 l 11,-5 6,-6 6,-17 v -12 l -6,-17 -11,-11 -17,-6 h -18 l -17,6 -5,6 -6,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12414" />
        <path
           d="m 3380,2676 v 120 l -57,-80 h 86"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12416" />
        <path
           d="m 3443,2768 v 5 l 6,12 6,5 11,6 h 23 l 11,-6 6,-5 6,-12 v -11 l -6,-12 -11,-17 -58,-57 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12418" />
        <path
           d="m 3626,2756 -6,-17 -11,-11 -17,-6 h -6 l -17,6 -12,11 -5,17 v 6 l 5,17 12,11 17,6 h 6 l 17,-6 11,-11 6,-23 v -28 l -6,-29 -11,-17 -17,-6 h -12 l -17,6 -6,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12420" />
        <path
           d="m 3666,2796 h 80 l -57,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12422" />
        <path
           d="m 3780,2728 h 103"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12424" />
        <path
           d="m 4003,2756 -6,-17 -11,-11 -17,-6 h -6 l -17,6 -11,11 -6,17 v 6 l 6,17 11,11 17,6 h 6 l 17,-6 11,-11 6,-23 v -28 l -6,-29 -11,-17 -17,-6 h -12 l -17,6 -5,11"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12426" />
        <path
           d="m 4043,2728 h 103"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12428" />
        <path
           d="m 4192,2676 v 120 h 40 l 17,-6 11,-11 6,-11 6,-18 v -28 l -6,-17 -6,-12 -11,-11 -17,-6 h -40"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12430" />
        <path
           d="m 4317,2688 -5,-6 5,-6 6,6"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12432" />
        <path
           d="m 4477,2676 v 120 l 46,-120 46,120 v -120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12434" />
        <path
           d="m 4615,2676 45,120 46,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12436" />
        <path
           d="m 4632,2716 h 57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12438" />
        <path
           d="m 4740,2676 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12440" />
        <path
           d="m 4786,2676 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12442" />
        <path
           d="M 4952,2796 V 2676"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12444" />
        <path
           d="m 4912,2796 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12446" />
        <path
           d="m 5015,2676 45,120 46,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12448" />
        <path
           d="m 5032,2716 h 57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12450" />
        <path
           d="m 5140,2676 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12452" />
        <path
           d="m 5186,2676 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12454" />
        <path
           d="m 1889,2453 46,120 45,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12456" />
        <path
           d="m 1906,2493 h 57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12458" />
        <path
           d="m 2123,2453 v 120 l 46,-120 46,120 v -120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12460" />
        <path
           d="m 2260,2453 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12462" />
        <path
           d="m 2306,2453 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12464" />
        <path
           d="m 2432,2453 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12466" />
        <path
           d="m 2478,2453 v 120 l 45,-120 46,120 v -120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12468" />
        <path
           d="m 2615,2573 v -85 l 5,-18 12,-11 17,-6 h 11 l 17,6 12,11 6,18 v 85"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12470" />
        <path
           d="m 2740,2453 v 120 l 46,-120 46,120 v -120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12472" />
        <path
           d="m 2986,2550 11,6 18,17 v -120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12474" />
        <path
           d="m 3083,2545 v 5 l 6,12 6,6 11,5 h 23 l 11,-5 6,-6 6,-12 v -11 l -6,-11 -11,-18 -58,-57 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12476" />
        <path
           d="m 3203,2590 -6,-5 -5,5 5,6 6,-6 v -11 l -6,-11 -5,-6"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12478" />
        <path
           d="m 3237,2590 -5,-5 -6,5 6,6 5,-6 v -11 l -5,-11 -6,-6"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12480" />
        <path
           d="m 3386,2573 46,-120 45,120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12482" />
        <path
           d="m 3500,2453 v 120 h 75"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12484" />
        <path
           d="m 3500,2516 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12486" />
        <path
           d="m 3500,2453 h 75"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12488" />
        <path
           d="m 3609,2453 v 120 h 51 l 17,-5 6,-6 6,-12 v -11 l -6,-11 -6,-6 -17,-6 h -51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12490" />
        <path
           d="m 3649,2516 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12492" />
        <path
           d="M 3769,2573 V 2453"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12494" />
        <path
           d="m 3729,2573 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12496" />
        <path
           d="m 3832,2453 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12498" />
        <path
           d="m 3963,2545 -6,11 -11,12 -11,5 h -23 l -12,-5 -11,-12 -6,-11 -6,-17 v -29 l 6,-17 6,-12 11,-11 12,-6 h 23 l 11,6 11,11 6,12"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12500" />
        <path
           d="m 3997,2453 46,120 46,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12502" />
        <path
           d="m 4015,2493 h 57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12504" />
        <path
           d="m 4123,2573 v -120 h 69"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12506" />
        <path
           d="m 4415,2545 -6,11 -12,12 -11,5 h -23 l -11,-5 -12,-12 -5,-11 -6,-17 v -29 l 6,-17 5,-12 12,-11 11,-6 h 23 l 11,6 12,11 6,12"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12508" />
        <path
           d="m 4449,2573 v -120 h 68"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12510" />
        <path
           d="m 4546,2453 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12512" />
        <path
           d="m 4546,2516 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12514" />
        <path
           d="m 4546,2453 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12516" />
        <path
           d="m 4655,2453 45,120 46,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12518" />
        <path
           d="m 4672,2493 h 57"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12520" />
        <path
           d="m 4780,2453 v 120 h 52 l 17,-5 6,-6 5,-12 v -11 l -5,-11 -6,-6 -17,-6 h -52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12522" />
        <path
           d="m 4820,2516 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12524" />
        <path
           d="m 4900,2453 46,120 46,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12526" />
        <path
           d="m 4917,2493 h 58"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12528" />
        <path
           d="m 5026,2453 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12530" />
        <path
           d="m 5237,2545 -5,11 -12,12 -11,5 h -23 l -11,-5 -12,-12 -6,-11 -5,-17 v -29 l 5,-17 6,-12 12,-11 11,-6 h 23 l 11,6 12,11 5,12"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12532" />
        <path
           d="m 5272,2453 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12534" />
        <path
           d="m 5272,2516 h 45"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12536" />
        <path
           d="m 5272,2453 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12538" />
        <path
           d="m 1889,2253 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12540" />
        <path
           d="m 1889,2316 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12542" />
        <path
           d="m 1992,2253 v 120 h 51 l 17,-5 6,-6 6,-12 v -11 l -6,-11 -6,-6 -17,-6 h -51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12544" />
        <path
           d="m 2032,2316 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12546" />
        <path
           d="m 2146,2373 -11,-5 -12,-12 -5,-11 -6,-17 v -29 l 6,-17 5,-12 12,-11 11,-6 h 23 l 11,6 12,11 6,12 5,17 v 29 l -5,17 -6,11 -12,12 -11,5 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12548" />
        <path
           d="m 2238,2253 v 120 l 45,-120 46,120 v -120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12550" />
        <path
           d="m 2535,2316 17,-6 6,-5 5,-12 v -17 l -5,-11 -6,-6 -17,-6 h -52 v 120 h 52 l 17,-5 6,-6 5,-12 v -11 l -5,-11 -6,-6 -17,-6 h -52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12552" />
        <path
           d="m 2637,2373 -11,-5 -11,-12 -6,-11 -6,-17 v -29 l 6,-17 6,-12 11,-11 11,-6 h 23 l 12,6 11,11 6,12 6,17 v 29 l -6,17 -6,11 -11,12 -12,5 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12554" />
        <path
           d="M 2769,2373 V 2253"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12556" />
        <path
           d="m 2729,2373 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12558" />
        <path
           d="M 2872,2373 V 2253"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12560" />
        <path
           d="m 2832,2373 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12562" />
        <path
           d="m 2969,2373 -12,-5 -11,-12 -6,-11 -5,-17 v -29 l 5,-17 6,-12 11,-11 12,-6 h 23 l 11,6 12,11 5,12 6,17 v 29 l -6,17 -5,11 -12,12 -11,5 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12564" />
        <path
           d="m 3060,2253 v 120 l 46,-120 46,120 v -120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12566" />
        <path
           d="m 3340,2373 -11,-5 -12,-12 -5,-11 -6,-17 v -29 l 6,-17 5,-12 12,-11 11,-6 h 23 l 12,6 11,11 6,12 5,17 v 29 l -5,17 -6,11 -11,12 -12,5 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12568" />
        <path
           d="m 3432,2253 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12570" />
        <path
           d="m 3432,2316 h 45"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12572" />
        <path
           d="m 3643,2253 v 120 h 52 l 17,-5 5,-6 6,-12 v -17 l -6,-11 -5,-6 -17,-6 h -52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12574" />
        <path
           d="m 3763,2253 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12576" />
        <path
           d="m 3809,2253 v 120 h 51 l 17,-5 6,-6 6,-12 v -17 l -6,-11 -6,-6 -17,-6 h -51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12578" />
        <path
           d="m 3929,2253 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12580" />
        <path
           d="m 3929,2316 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12582" />
        <path
           d="m 3929,2253 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12584" />
        <path
           d="m 4049,2259 -6,-6 -6,6 6,6 6,-6 v -11 l -6,-12 -6,-6"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12586" />
        <path
           d="m 4203,2373 29,-120 28,120 29,-120 28,120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12588" />
        <path
           d="m 4340,2253 46,120 46,-120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12590" />
        <path
           d="m 4357,2293 h 58"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12592" />
        <path
           d="M 4506,2373 V 2253"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12594" />
        <path
           d="m 4466,2373 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12596" />
        <path
           d="m 4569,2253 v 120 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12598" />
        <path
           d="m 4569,2316 h 46"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12600" />
        <path
           d="m 4569,2253 h 74"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12602" />
        <path
           d="m 4677,2253 v 120 h 52 l 17,-5 6,-6 5,-12 v -11 l -5,-11 -6,-6 -17,-6 h -52"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12604" />
        <path
           d="m 4717,2316 40,-63"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12606" />
        <path
           d="m 4940,2373 -11,-5 -12,-12 -5,-11 -6,-17 v -29 l 6,-17 5,-12 12,-11 11,-6 h 23 l 12,6 11,11 6,12 5,17 v 29 l -5,17 -6,11 -11,12 -12,5 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12608" />
        <path
           d="m 5032,2253 v 120 l 80,-120 v 120"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12610" />
        <path
           d="M 1929,2173 V 2053"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12612" />
        <path
           d="m 1889,2173 h 80"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12614" />
        <path
           d="m 2026,2173 -11,-5 -12,-12 -5,-11 -6,-17 v -29 l 6,-17 5,-12 12,-11 11,-6 h 23 l 11,6 12,11 6,12 5,17 v 29 l -5,17 -6,11 -12,12 -11,5 h -23"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12616" />
        <path
           d="m 2118,2053 v 120 h 51 l 17,-5 6,-6 6,-12 v -17 l -6,-11 -6,-6 -17,-6 h -51"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12618" />
        <path
           d="M 624,4019 H 5501"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12620" />
        <path
           d="M 624,3555 H 5501"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12622" />
        <path
           d="M 624,3091 H 5501"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12624" />
        <path
           d="M 624,4019 V 1981 h 4877"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12626" />
        <path
           d="M 1817,3555 V 1981"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12628" />
        <path
           d="M 5501,4019 V 1981"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12630" />
        <g
           id="g12632">
          <path
             d="m 1261,15671 -88,-46 298,-354 z m -88,-46 298,-354 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12634" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46487,-0.88538,-0.88538,-0.46487,1179,15616)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#139b48;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12638"><tspan
             x="0 74.565788 149.13158 174.7468 212.02969 301.48181"
             y="0"
             sodipodi:role="line"
             id="tspan12636">20' SW</tspan></text>
        <g
           id="g12640">
          <path
             d="m 3348,8531 -87,-47 203,-174 z m -87,-47 203,-174 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12642" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46402,-0.88582,-0.88582,-0.46402,3257,8494)"
           style="font-variant:normal;font-weight:normal;font-size:134.11px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00bfff;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12646"><tspan
             x="0 96.827736 134.11044"
             y="0"
             sodipodi:role="line"
             id="tspan12644">R/W</tspan></text>
        <g
           id="g12648">
          <path
             d="m 3583,10367 45,-85 65,142 z m 45,-85 65,142 44,-85 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12650" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88475,0.46606,0.46606,-0.88475,3627,10281)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12654"><tspan
             x="0"
             y="0"
             id="tspan12652">W</tspan></text>
        <g
           id="g12656">
          <path
             d="m 7667,5637 -88,-46 298,-353 z m -88,-46 298,-353 -88,-47 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12658" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46487,-0.88538,-0.88538,-0.46487,7585,5582)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#139b48;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12662"><tspan
             x="0 74.565788 149.13158 174.7468 212.02969 301.48181"
             y="0"
             sodipodi:role="line"
             id="tspan12660">20' SW</tspan></text>
        <g
           id="g12664">
          <path
             d="m 3215,13262 v -648 l 3575,648 z m 0,-648 3575,648 v -648 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12666" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,3267,13080)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12670"><tspan
             x="0 121.03464 251.457 372.49164 493.52628 605.34082 726.37543 828.80225 875.40564 996.44025 1126.8627 1247.8972 1368.9319 1489.9666 1536.5699 1638.9967 1685.6001 1788.0269 1918.4492 1965.0526 2076.8672 2188.6816 2235.2852 2347.0996 2449.5264 2496.1299 2617.1646"
             y="0"
             sodipodi:role="line"
             id="tspan12668">CONNECT CONDUIT TO EXISTING</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,3273,12878)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12674"><tspan
             x="0 93.206726 152.71822 199.32158 255.14503 366.95959 487.99423 534.5976 646.41211 758.22668 860.6535 972.46802 1028.2915 1074.8949 1186.7094 1298.5239 1419.5586 1466.162 1577.9764 1689.791 1848.0413 1959.8558 2080.8904 2127.4939 2220.7007 2332.5151 2434.9419 2546.7566 2667.791 2779.6057"
             y="0"
             sodipodi:role="line"
             id="tspan12672">4&quot; (PRIVATE) PVC SEWER LATERAL</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,3262,12676)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12678"><tspan
             x="0 121.03464 232.84918 335.276 447.09055 568.12518 679.93976 800.97437 922.00897 1033.8235 1080.4269 1192.2415 1331.8839 1452.9186 1564.733 1611.3364 1704.5432 1751.1466 1862.9611 1993.3834 2114.4182 2170.2415 2263.4482 2356.655 2449.8618 2543.0684 2636.2751 2729.4819"
             y="0"
             sodipodi:role="line"
             id="tspan12676">REFERENCE EMRA # AGR-0000874</tspan></text>
        <g
           id="g12680">
          <path
             d="m 1846,13358 -105,61 119,-24 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12682" />
        </g>
        <path
           d="m 1853,13377 1151,-439 h 163"
           style="fill:none;stroke:#000000;stroke-width:17;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12684" />
        <g
           id="g12686">
          <path
             d="m 5715,10707 v -278 l 2452,278 z m 0,-278 2452,278 v -278 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12688" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,5765,10525)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12692"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12690">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,6063,10525)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12696"><tspan
             x="0 93.206726 152.71822 199.32158 311.13614 422.95068 543.98529 655.79987 758.22668 851.43341 981.85577 1140.1061 1186.7094 1326.3518 1438.1664 1559.201 1605.8044 1708.2312 1838.6536 1931.8604"
             y="0"
             sodipodi:role="line"
             id="tspan12694">1&quot; BACKFLOW MANIFOLD</tspan></text>
        <g
           id="g12698">
          <path
             d="m 4559,10608 -118,28 121,12 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12700" />
        </g>
        <path
           d="m 4561,10628 942,-60 h 164"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12702" />
        <g
           id="g12704">
          <path
             d="m 5976,11058 v -277 l 1661,277 z m 0,-277 1661,277 v -277 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12706" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,6026,10876)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12710"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12708">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,6340,10876)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12714"><tspan
             x="0 158.25027 270.06482 372.49164 484.30618 605.34082 651.94415 791.58661 903.40118 1005.828 1117.6426"
             y="0"
             sodipodi:role="line"
             id="tspan12712">WATER METER</tspan></text>
        <g
           id="g12716">
          <path
             d="m 5243,10969 -116,36 122,4 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12718" />
        </g>
        <path
           d="m 5246,10989 518,-70 h 164"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12720" />
        <g
           id="g12722">
          <path
             d="m 596,9205 v -277 l 2158,277 z m 0,-277 2158,277 v -277 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12724" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,646,9023)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12728"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12726">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,962,9023)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12732"><tspan
             x="0 111.81454 232.84918 353.88382 474.91846 605.34082 726.37543 838.19 959.22461 1005.828 1117.6426 1229.457 1341.2716 1443.6985 1490.3019 1611.3364"
             y="0"
             sodipodi:role="line"
             id="tspan12730">ANCHORED SEATING</tspan></text>
        <path
           d="m 3184,9028 -219,39 h -163"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12734" />
        <g
           id="g12736">
          <path
             d="m 922,9964 v -447 l 1377,447 z m 0,-447 1377,447 v -447 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12738" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,972,9782)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12742"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12740">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1288,9782)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12746"><tspan
             x="0 111.81454 232.84918 353.88382 474.91846 605.34082 726.37543 838.19"
             y="0"
             sodipodi:role="line"
             id="tspan12744">ANCHORED</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1513,9579)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12750"><tspan
             x="0 111.81454 223.62909 335.44363 437.87045 484.47382 605.50848"
             y="0"
             sodipodi:role="line"
             id="tspan12748">SEATING</tspan></text>
        <g
           id="g12752">
          <path
             d="m 2666,9836 115,-40 -122,1 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12754" />
        </g>
        <path
           d="m 2662,9817 -152,26 h -163"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12756" />
        <g
           id="g12758">
          <path
             d="m 591,9459 v -278 l 1954,278 z m 0,-278 1954,278 v -278 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12760" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,641,9276)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12764"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12762">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,957,9276)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12768"><tspan
             x="0 111.81454 232.84918 353.88382 474.91846 605.34082 726.37543 838.19 959.22461 1005.828 1108.2548 1220.0693 1331.8839 1425.0907"
             y="0"
             sodipodi:role="line"
             id="tspan12766">ANCHORED TABLE</tspan></text>
        <path
           d="m 2938,9380 -181,-59 h -164"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12770" />
        <g
           id="g12772">
          <path
             d="m 1482,8971 v -278 l 1184,278 z m 0,-278 1184,278 v -278 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12774" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1531,8789)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12778"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12776">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1835,8789)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12782"><tspan
             x="0 111.81454 205.02127 316.83582 437.87045 540.2973 652.11182"
             y="0"
             sodipodi:role="line"
             id="tspan12780">PLANTER</tspan></text>
        <g
           id="g12784">
          <path
             d="m 3114,8807 114,-43 -122,4 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12786" />
        </g>
        <path
           d="m 3110,8787 -232,46 h -164"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12788" />
        <g
           id="g12790">
          <path
             d="m 982,8063 v -278 l 2006,278 z m 0,-278 2006,278 v -278 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12792" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1032,7880)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12796"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12794">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1349,7880)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12800"><tspan
             x="0 111.81454 232.84918 353.88382 474.91846 605.34082 726.37543 838.19 959.22461 1005.828 1117.6426 1229.457 1350.4917 1471.5264"
             y="0"
             sodipodi:role="line"
             id="tspan12798">ANCHORED BENCH</tspan></text>
        <g
           id="g12802">
          <path
             d="m 3456,8118 112,50 -89,-83 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12804" />
        </g>
        <path
           d="M 3468,8102 3200,7925 H 3036"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12806" />
        <g
           id="g12808">
          <path
             d="m 4759,11979 v -649 l 3998,649 z m 0,-649 3998,649 v -649 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12810" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,4806,11797)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12814"><tspan
             x="0 111.81454 232.84918 363.27155 475.08609 605.50848 717.323 829.13757 950.17218 996.77557 1089.9823 1183.189 1215.2079 1261.8113 1364.238 1485.2727 1597.0873 1718.1218 1839.1565"
             y="0"
             sodipodi:role="line"
             id="tspan12812">PROPOSED 50' TRENCH</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,4815,11594)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12818"><tspan
             x="0 102.42682 232.84918 279.45255 391.26709 484.47382 596.28839 717.323 829.13757 875.74091 968.94763 1028.4591 1075.0625 1130.886 1242.7004 1363.7351 1410.3385 1522.1531 1633.9675 1736.3944 1848.209 1904.0323 1950.6357 2062.4502 2174.2649 2295.2996 2341.9028 2453.7173 2565.532 2723.7822 2835.5967 2956.6313 3003.2349 3096.4414 3208.2561 3310.6829 3422.4973 3543.532 3655.3467"
             y="0"
             sodipodi:role="line"
             id="tspan12816">TO PLACE 4&quot; (PRIVATE) PVC SEWER LATERAL</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,4805,11392)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12822"><tspan
             x="0 121.03464 232.84918 335.276 447.09055 568.12518 679.93976 800.97437 922.00897 1033.8235 1080.4269 1192.2415 1331.8839 1452.9186 1564.733 1611.3364 1704.5432 1751.1466 1862.9611 1993.3834 2114.4182 2170.2415 2263.4482 2356.655 2449.8618 2543.0684 2636.2751 2729.4819"
             y="0"
             sodipodi:role="line"
             id="tspan12820">REFERENCE EMRA # AGR-0000874</tspan></text>
        <g
           id="g12824">
          <path
             d="m 3227,10849 -113,-43 93,78 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12826" />
        </g>
        <path
           d="m 3217,10867 1330,787 h 164"
           style="fill:none;stroke:#000000;stroke-width:17;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12828" />
        <g
           id="g12830">
          <path
             d="m 7842,12606 46,-88 1127,704 z m 46,-88 1127,704 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12832" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.8852,0.46521,0.46521,-0.8852,7891,12521)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12836"><tspan
             x="0 89.452011 178.90402 216.18686 305.63889 387.58066 424.86353 521.69165 626.02997 663.31281 737.87848 785.48792 822.77075 949.37146 1038.8235 1120.7653 1210.2173"
             y="0"
             sodipodi:role="line"
             id="tspan12834">EXISTING 1&quot; WATER</tspan></text>
        <g
           id="g12838">
          <path
             d="m 7516,7287 -88,-46 216,-198 z m -88,-46 216,-198 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12840" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46776,-0.88386,-0.88386,-0.46776,7427,7247)"
           style="font-variant:normal;font-weight:normal;font-size:134.112px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12844"><tspan
             x="0 96.828522 186.28091"
             y="0"
             sodipodi:role="line"
             id="tspan12842">C&amp;G</tspan></text>
        <g
           id="g12846">
          <path
             d="m 6914,9912 v -278 l 987,278 z m 0,-278 987,278 v -278 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12848" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,6964,9730)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12852"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12850">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,7268,9730)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12856"><tspan
             x="0 111.81454 223.62909 344.66373 465.69836"
             y="0"
             sodipodi:role="line"
             id="tspan12854">BENCH</tspan></text>
        <g
           id="g12858">
          <path
             d="m 5413,8926 -112,-48 91,81 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12860" />
        </g>
        <path
           d="m 5402,8943 1300,830 h 164"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12862" />
        <g
           id="g12864">
          <path
             d="m 7740,8183 v -277 l 988,277 z m 0,-277 988,277 v -277 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12866" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,7790,8001)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12870"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12868">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,8094,8001)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12874"><tspan
             x="0 111.81454 223.62909 344.66373 465.69836"
             y="0"
             sodipodi:role="line"
             id="tspan12872">BENCH</tspan></text>
        <g
           id="g12876">
          <path
             d="m 6277,7280 -113,-44 93,78 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12878" />
        </g>
        <path
           d="m 6267,7297 1262,747 h 163"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12880" />
        <g
           id="g12882">
          <path
             d="m 2150,5944 v -278 l 2005,278 z m 0,-278 2005,278 v -278 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12884" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,2200,5761)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12888"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12886">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,2516,5761)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12892"><tspan
             x="0 111.81454 232.84918 353.88382 474.91846 605.34082 726.37543 838.19 959.22461 1005.828 1117.6426 1229.457 1350.4917 1471.5264"
             y="0"
             sodipodi:role="line"
             id="tspan12890">ANCHORED BENCH</tspan></text>
        <g
           id="g12894">
          <path
             d="m 4578,5973 110,51 -88,-84 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12896" />
        </g>
        <path
           d="M 4589,5957 4367,5806 H 4203"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12898" />
        <g
           id="g12900">
          <path
             d="m 1946,6293 v -277 l 1952,277 z m 0,-277 1952,277 v -277 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12902" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1996,6111)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12906"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12904">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,2313,6111)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12910"><tspan
             x="0 111.81454 232.84918 353.88382 474.91846 605.34082 726.37543 838.19 959.22461 1005.828 1126.8627 1247.8972 1359.7118 1406.3152"
             y="0"
             sodipodi:role="line"
             id="tspan12908">ANCHORED CHAIR</tspan></text>
        <g
           id="g12912">
          <path
             d="m 4154,6895 30,118 10,-121 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12914" />
        </g>
        <path
           d="m 4174,6894 -64,-738 h -164"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12916" />
        <g
           id="g12918">
          <path
             d="m 3657,13947 v -277 l 860,277 z m 0,-277 860,277 v -277 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12920" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,3707,13765)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12924"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan12922">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,4019,13765)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12928"><tspan
             x="0 102.42682 223.46146 335.276"
             y="0"
             sodipodi:role="line"
             id="tspan12926">TREE</tspan></text>
        <g
           id="g12930">
          <path
             d="m 2494,14204 -102,66 118,-30 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12932" />
        </g>
        <path
           d="m 2502,14222 943,-413 h 164"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12934" />
        <g
           id="g12936">
          <path
             d="M 576,7505 V 6457 l 2922,1048 z m 0,-1048 2922,1048 V 6457 Z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12938" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,712,7323)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12942"><tspan
             x="0 55.823456 176.85809 232.68155 279.28491 335.10837 446.92291 567.95752 614.56091 726.37543 838.19 940.61682 1052.4314 1108.2548 1154.8582 1266.6727 1378.4873 1536.7375 1648.5521 1769.5867 1816.1901 1937.2247 2030.4314 2142.2461 2254.0605 2375.0952 2505.5176 2626.5522"
             y="0"
             sodipodi:role="line"
             id="tspan12940">(N) (PRIVATE) SEWER CLEANOUT</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1705,7121)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12946"><tspan
             x="0 111.81454 223.62909 344.66373 391.26709 512.30176 558.90509 661.33191 773.14648 819.74982 931.56439 1033.9912 1145.8058 1266.8403 1387.875 1499.6896 1620.7242"
             y="0"
             sodipodi:role="line"
             id="tspan12944">PER CITY STANDARD</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1992,6919)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12950"><tspan
             x="0 111.81454 232.84918 344.66373 400.48718 493.69391 586.90063 680.10736 726.71075 773.31409 885.12866 1006.1633 1117.9778 1173.8013 1267.0081 1360.2147"
             y="0"
             sodipodi:role="line"
             id="tspan12948">SDS-101, SDS-103</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,623,6717)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12954"><tspan
             x="0 121.03464 232.84918 335.276 447.09055 568.12518 679.93976 800.97437 922.00897 1033.8235 1080.4269 1192.2415 1331.8839 1452.9186 1564.733 1611.3364 1704.5432 1751.1466 1862.9611 1993.3834 2114.4182 2170.2415 2263.4482 2356.655 2449.8618 2543.0684 2636.2751 2729.4819"
             y="0"
             sodipodi:role="line"
             id="tspan12952">REFERENCE EMRA # AGR-0000874</tspan></text>
        <g
           id="g12956">
          <path
             d="m 4091,7441 121,-9 -117,-31 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12958" />
        </g>
        <path
           d="m 4093,7421 -384,-36"
           style="fill:none;stroke:#000000;stroke-width:17;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12960" />
        <g
           id="g12962">
          <path
             d="m 4354,8112 96,75 -67,-102 z"
             style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12964" />
        </g>
        <path
           d="M 4369,8099 3709,7385 H 3546"
           style="fill:none;stroke:#000000;stroke-width:17;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path12966" />
        <g
           id="g12968">
          <path
             d="m 1490,12068 -88,-46 204,-174 z m -88,-46 204,-174 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12970" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46699,-0.88426,-0.88426,-0.46699,1399,12032)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00bfff;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12974"><tspan
             x="0 96.827919 134.11069"
             y="0"
             sodipodi:role="line"
             id="tspan12972">R/W</tspan></text>
        <g
           id="g12976">
          <path
             d="M 7009,9511 V 8459 l 4991,1052 z m 0,-1052 4991,1052 V 8459 Z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path12978" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,7056,9329)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12982"><tspan
             x="0 121.03464 232.84918 372.49164 502.914 614.72852 726.54309 773.14648 884.961 1005.9957 1127.0303 1173.6337 1294.6683 1406.4828 1518.2974 1611.5042 1723.3186 1844.3533 1956.1678 2002.7712 2095.978 2189.1846 2282.3914 2328.9946 2440.8093 2571.2317 2673.6584 2776.0852 2822.6887 2934.5032 2981.1064 3102.1411 3213.9558 3372.2061 3484.0205 3577.2273 3689.0417 3735.6453 3847.4597 3959.2742 4080.3088 4192.1235 4285.3301"
             y="0"
             sodipodi:role="line"
             id="tspan12980">REMOVE AND REPLACE 915 SQFT SIDEWALK PANEL,</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,7115.6034,9127)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12986"><tspan
             x="0 111.81454 158.41791 279.45255 391.26709 549.51733 661.33191 754.53864 866.35321 912.95654 1052.599 1173.6337 1285.4482 1387.875 1434.4784 1546.293 1658.1074 1704.7108 1825.7455 1937.5601 2049.3745 2161.1892 2207.7925 2328.8271 2440.6416 2561.6763 2608.2795 2729.3142 2841.1289 2952.9434 3046.1501 3157.9646 3278.9993 3390.8137 3511.8484 3558.4519 3642.2708 3772.6931 3819.2966 3940.3313 4042.7581 4089.3613 4191.7881"
             y="0"
             sodipodi:role="line"
             id="tspan12984">SIDEWALK MUST BE REPAIRED/REPLACED JOINT TO</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,7065,8925)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12990"><tspan
             x="0 83.819 214.24136 260.84473 381.87936 484.30618 530.90955 577.51294 689.32745 801.14203 922.17664 1033.9912 1127.1979 1239.0125 1285.6158 1425.2583 1546.293 1658.1074 1760.5343 1807.1377 1918.9521 2030.7667 2077.3701 2179.7969 2273.0037 2394.0383 2505.8528 2626.8875 2673.4907 2831.7412 2878.3445 2980.7712 3101.8059 3148.4092 3260.2239 3381.2585 3502.2932 3623.3276 3753.75 3874.7847 3995.8193 4116.854 4163.4575 4284.4922"
             y="0"
             sodipodi:role="line"
             id="tspan12988">JOINT. PANELS MUST BE FLUSH WITH SURROUNDING</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,7062,8723)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12994"><tspan
             x="0 111.81454 158.41791 279.45255 391.26709 549.51733 661.33191 754.53864 866.35321 912.95654 1024.7711 1145.8058 1266.8403 1313.4437 1443.8661 1564.9008 1676.7153 1723.3186 1835.1332 1956.1678 2086.5901 2189.0171 2310.0518 2421.8662 2542.9009 2589.5042 2636.1077 2775.75 2887.5645 2934.168 3055.2026 3157.6294 3269.4438 3316.0474 3437.082 3483.6853 3595.4998 3716.5344 3846.9568 3967.9915 4014.5947 4135.6294"
             y="0"
             sodipodi:role="line"
             id="tspan12992">SIDEWALK AND ONE ANOTHER. MAINTAIN SCORING</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,7056,8521)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text12998"><tspan
             x="0 111.81454 223.62909 326.05591 428.48273 540.2973 661.33191 782.36652 828.96991 959.39227 1061.8191 1108.4225 1220.2371 1332.0515 1378.6549 1490.4695 1592.8962 1639.4996 1760.5343 1890.9567 1937.5601 2049.3745 2170.4092 2291.4438 2412.4785 2542.9009 2663.9355 2784.9702 2906.0046 2952.6082 3073.6428 3204.0652 3250.6685 3362.4829 3409.0864 3530.1211 3641.9355 3800.1858 3912.0005 4005.207"
             y="0"
             sodipodi:role="line"
             id="tspan12996">PATTERN OF EXISTING SURROUNDING SIDEWALK</tspan></text>
        <path
           d="m 5434,8081 -27,-167"
           style="fill:none;stroke:#000000;stroke-width:17;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13000" />
        <path
           d="m 5421,7997 1377,988 h 163"
           style="fill:none;stroke:#000000;stroke-width:17;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13002" />
        <path
           d="m 699,4631 v -447 h 3751 v 447 H 699"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13004" />
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,751,4449)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13008"><tspan
             x="0 130.42236 251.457 344.66373 456.47827 503.08163 661.33191 791.75427 912.78894 1024.6035 1071.2068 1117.8102 1238.8448 1285.4482 1387.875 1508.9097 1620.7242 1667.3275 1779.1421 1900.1768 2011.9913 2105.198 2151.8013 2272.8359 2319.4395 2440.4741 2487.0774 2617.4998 2738.5344 2840.9612 2887.5645 3017.9868 3120.4138 3167.0171 3325.2673 3437.082"
             y="0"
             sodipodi:role="line"
             id="tspan13006">ONLY WORK IN THE PUBLIC RIGHT OF WAY</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,747,4247)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13012"><tspan
             x="0 139.64246 251.457 363.27155 409.87491 521.68945 633.50403 680.10736 791.92194 903.73645 1024.7711 1127.1979 1257.6202 1378.6549 1518.2974 1630.1119 1751.1466 1797.7499 1928.1722 2049.207 2095.8103 2198.2371 2319.2717 2365.875 2477.6897 2524.293 2636.1077 2747.9221 2868.9568 3008.5991 3055.2026"
             y="0"
             sodipodi:role="line"
             id="tspan13010">MAY BE PERFORMED ON THIS PERMIT</tspan></text>
        <g
           id="g13014">
          <path
             d="m 7710,17565 -88,-46 132,-39 z m -88,-46 132,-39 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13016" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46062,-0.8876,-0.8876,-0.46062,7625,17516)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13020"><tspan
             x="0"
             y="0"
             id="tspan13018">S</tspan></text>
        <g
           id="g13022">
          <path
             d="m 2978,14218 121,-231 1691,1183 z m 121,-231 1691,1183 121,-231 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13024" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88533,0.46496,0.46496,-0.88533,3131,14188)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13028"><tspan
             x="0 89.451904 178.90381 216.18661 305.63852 387.5802 424.86301 521.69104 626.02924 663.31201 737.87762 785.48694 822.76978 867.42865 956.88055 1053.7085 1090.9913 1180.4432 1269.8951 1351.8369 1441.2888 1485.9476 1523.2305 1612.6824 1702.1343"
             y="0"
             sodipodi:role="line"
             id="tspan13026">EXISTING 4&quot; (PRIVATE) PVC</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(0.88538,0.46487,0.46487,-0.88538,3506,14202)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13032"><tspan
             x="0 89.452118 178.90424 305.50516 394.95728 491.78549 529.06836 603.63416 693.0863 775.0282 864.48029 961.30853 1050.7606"
             y="0"
             sodipodi:role="line"
             id="tspan13030">SEWER LATERAL</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1303,10509)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13036"><tspan
             x="0 93.206726 186.41345 279.62018"
             y="0"
             sodipodi:role="line"
             id="tspan13034">5636</tspan></text>
        <path
           d="m 1752,10604 v -156 h -492"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13038" />
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1005,7060)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13042"><tspan
             x="0 93.206726 186.41345 279.62018"
             y="0"
             sodipodi:role="line"
             id="tspan13040">5630</tspan></text>
        <path
           d="M 1454,7155 V 6999 H 961"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13044" />
        <path
           d="m 718,5171 v -446 h 2249 v 446 H 718"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13046" />
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,1053,4989)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13050"><tspan
             x="0 121.03464 232.84918 335.276 447.09055 568.12518 679.93976 800.97437 922.00897 1033.8235 1080.4269 1192.2415 1331.8839 1452.9186"
             y="0"
             sodipodi:role="line"
             id="tspan13048">REFERENCE EMRA</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,918,4787)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13054"><tspan
             x="0 121.03464 242.06927 381.71173 493.52628 605.34082 726.37543 772.97882 884.79333 1015.2157 1136.2504 1192.0739 1285.2805 1378.4873 1471.694 1564.9008 1658.1074 1751.3142"
             y="0"
             sodipodi:role="line"
             id="tspan13052">NUMBER AGR-0000874</tspan></text>
        <g
           id="g13056">
          <path
             d="m 9079,11954 h -277 l 416,-239 z m -277,0 416,-239 h -554 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13058" />
        </g>
        <g
           id="g13060">
          <path
             d="m 9218,11715 h -554 l 415,-240 z m -554,0 415,-240 h -277 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13062" />
        </g>
        <path
           d="m 8802,11954 -138,-239 138,-240 h 277 l 139,240 -139,239 h -277"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13064" />
        <path
           d="m 8664,11715 h 554"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13066" />
        <path
           d="m 8941,11715 v 239"
           style="fill:none;stroke:#000000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13068" />
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,8809,11773)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13072"><tspan
             x="0"
             y="0"
             id="tspan13070">1</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,8987,11773)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13076"><tspan
             x="0 74.56572"
             y="0"
             sodipodi:role="line"
             id="tspan13074">4&quot;</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,8878,11554)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13080"><tspan
             x="0 74.56572 149.13144"
             y="0"
             sodipodi:role="line"
             id="tspan13078">50'</tspan></text>
      </g>
    </g>
    <g
       id="g13082">
      <g
         id="g13084"
         clip-path="url(#clipPath13088)" />
    </g>
    <g
       id="g13090">
      <g
         id="g13092"
         clip-path="url(#clipPath13096)">
        <g
           id="g13098"
           transform="matrix(122,0,0,121,3366,10155)">
          <image
             width="1"
             height="1"
             style="image-rendering:optimizeSpeed"
             preserveAspectRatio="none"
             transform="matrix(1,0,0,-1,0,1)"
             xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAACkAAAApCAYAAACoYAD2AAAABHNCSVQICAgIfAhkiAAADKlJREFUWIWtmdmvbcdRxn/V3WvY8zn3jNfXw7WvnWCSyCSyAhb8LxEvICI5xvGAHERwEozkRIIIJAQPIKQ8IZAQbzxZQgIlGAFRjJ3E8x18fXzOPtOe11rdXTz02ufeEB6QTUlLe9Daq7+uqq/qq97CdqZMGsqYkXkAJRCpiFAKMSoaADXQ34KQw+4+RAPdHcoX/ohK+qgoELEasTSUvqYbVhx84+sQKphPIBM4HtMvHX55zICAoWbJiomLMCKZAgKcQ+FB6KAo2BVsZT0yazldTbCjIdP5BIxDNrbQ0wqyLgx3+OKzzzPZ3uZmbQnlvVTSQyWCRETBqsdpQydUdOoln9reIBzcpLp5nVe/99dweAChJrPCto2crg5ZlU0CVrZAV0AFRQShQAmwXfSp5jMEyLs9xlUF/QEEB9kQfMkTX3kGs72L7F3mtaPbDB64xngCjRREAZXWA0RAsVpjfUXRLAknRzx6ZZ94OqY6PuSNv/87ePdtWEzolobF8hhijRHajUJuoQkgZEY3Ni+xOhyTtZuYAVr0oBhCucXnn/46ndEVbH+Tn968Tb6zwXnmmcVIlm8QxLUgBcQkoJKAEmrKTgGrGYPcMvnoNqNOgfE1VwvhB7/7HKxmcHzEwIHUE2wb8bq9BOM0zy1mVWGBoltyUgXobMD2Vb7wtW8zy7d589Y5o+19Lu3vc3B6AIVCptR1TRSDYlqAAhgwJu24qqBwEBukW6DLBeIEnU7I6imfsSt++PzTIDky/og9KhwrkIyxrliJQTrdvq4WM3rWUcVIIxY6I9i5j3u/9CRnGw8QN++HcpvFypN3OtTjD2CzBOshVm14DeDaeLt0GRJoZyF6UIVqCZmBzNLNIu74HR7Wmv946nmyvCQb32BIjXGWQ3+GtwZxoP3+gLPZEooeSA6b+zz0G08z+twvc0t7HNUOyg1YVMlbXQe+guUplAHwif3qQO1d7wVrLaFpILQgMwtG0/s4Aztlg4rHouWfvvwkSCSbjfE6Jesaaj/FOOB8Nof+BkgXtq/y6d98jtGjj/Pm8YKl5DCbgF/CqIDVGRiBqobBCLB3PIeAgo2GPEARFJlXFEEY5D16RZeeK3HR4MRBVsJolzM34PVF4AvffAl6fRqXYzZ2qFc1KMgAdGZyNBtBuc2vvvznnPS2+PHBKZsPXeN0tbyLCOZOWDVL35kqeTKaBDAYXExArSamJouoxJZg6bWyoJkAgW5s2FlO2Zuf8OrvPQtxCfMjkHlaQkUg68Hla7zncz7QLr2HPsPpeAKAUGF1gdUJME9FTGMKazQQXRticweUxARePEiNGk80gWAbgm3wtkGNQm1xnV0WwXG9Chx3R7B7BYIB20G8wZjhEFwHigGf++rvcLuxNMNd5kcT2NjFaiSPFUWck+mcPK6wsUFiAyG2INMlMTFaBbyJ1C6yygKLPLDIAvPcs8o9VRHwRQAbKYs+/r0D9q48Ao3hmJyHf+spsF3oXMLQwXrNXqTo88S3vsP1kLMY7CMbO0TXgcUMK4GMCpEaEUWxiFqsZogatPW1qACa7hFQUbxRgoVoFLURbEwpvM4atYQZ9PobnB4fUmxfoiwyes7xyGOf59Yrr6DeYyhGcGmfuj+k6XTo723T3L4B4zHDnV2MGqJmeCmpTUEgI2IxEZwqRkE05ZtKilIwEGwiOhcF3qVrnc+aAQYlYmyE5YrgBa85N05m9K89Clt7UA4wZEN+5annuDVdUmeW2ds/przvCrKzyeT2AagjUlBJFy8dvClQXHKGpn6tJt5FrnVr5I7LtEUcMvDt1WQQMvJexnQyZnjfFfzpKV4sMtji+9dv8NCTvw39AY57HsQPtlAMNjP0Hr6X+fW36G3dzzLLiCheLJgGTEydLq5Zm1iKiRcMvlAxmLaFJzIZNYhKy3iDUfA2UjOl8+AOk9sfkm1vYYuSeX3A5kPXcHkDvR6GScP1RcB2RpRZl/mNm3S2RizmZ5Ap3hgwbYhilpgMBBMJxif183MA77yuAdpWNNhoUmrGthKUjuXkBDoZrnBM3n+H3j2XWYrw5o3b7Hzz20jxvddUgDyAqKA4KmuoXJbAiU0LBpAYyNSDNATjCUJbLw0/Zxf18U5ZMvqzn72NkLepEiNEhQguRoxGhIiL4KqiCyFiolKE5A1r2vyyMSVYTI7KY8TFSLCR2oREiqh3AfrfLBEKSJtae3ydsmrSd236CLElY2oajdhWBQgEiXiTdnnxGG27jLa80FQDNSmHdhXhY5u2mIWL/DURooDBgApBDG4dKi9gJbk+/syOPe1P7nr2Wun8P9h6GV1v17TYBRXTgmx1YJBIbSKGSFizVdswtB5VgagmbULNJ3IitK1f4x1wLQkjJmVBG2WXQKTPQQ1hPQZc5Elod5mARtMK3DYN0gbi/1z//2xrEaKSwKX11+o+3eOI8SLx70afLICm4cq0O02+NoC9SPaPa6bdvLQhDpKidZHqAqjHEer0C2nl/3oMIIJKCsma3uJQIipuvaP2iR8fKLTSDdcOcnfPSB4ImC0HebOE+YyizKFagW+4tLsP55O2HCQyxVYHJk+vVcLHtyjgsozKNxT9bipnYmA2AwnQLDHUGP/RTfZLx+XdTarDA+h3ISs5OTiCcnDRwmgJddFh9K7rE9h8MQOU+dkp2WiYxoytTfb392A1pVtPMed//DKMb6OTMfgVzkiaP1aezZ191vVQpZVld5FKPlmUUQHplJheD6yjqT3Mp1AvOfjJG8hyykYzxzAfc22jJFtN2d3daqc6AeNYzFYYdYC5E+a7jlMM8a7x4GOaEWKMmOEghXm0yXZ3AOMjfu1T17j1ja9h6DuOXv9PhrGiOjvCL5bYogApqM5XrVSz7VzdPljaM59Wqn0SU1XwHokKTU0WIkwm3Ls54sarP4DFFMNHt/ivv/wz9gY5fj7FWUGjQKNkvdGdEXVNEoltWVJMK3o/tglYayHLCIsFrjckzuYsDsc8uLnF9T/9EwgNDr+EJYxvvM/le36BcdHhzHsIARGbTifk57tLEgKfjN0AYVVDVgCWYdHBBmXk4OTd92BVQTVdq4vAj77zEozfZ3X2AWIbZDSkXi4xSgrrRS1MdTS2w1awsS2+DsiR6NpxNmC1QaQCaU/MjLlTB9e1tz2OKfKM84NbFLMz3PiA11/+A6AGX2GKKpDVEZoT3v7DZ7hnuERXB+j0GIoCpw1xNqG0ILmFRqAx1EapSwMZ4AyYAiixoUMWDE4rnMywcYK1VTqOKUrwClkOWkEWodsFsYg2XOlm7NXn/OSlFyBfwuIQWGCGxQbqFwypoBozmt+m05xw79XLcDZmo1Mw6Jes5lO0SSNsub0PeQH1MhVds5Z0DqM2jQqkjlEU7bFKloHJoDfC2RxiA5PTBLaa4BannL/3OsPVMegMVicQlqAegS21WUSaU8x+nzoUXH32ZXT4GPnoPsanR8xzqLc70OnBxMDJDHLDcLNg0pylUPs+hAznwVKhdkK0S3zwUPQh24RFhEUDcUW5adgcFpycHDMwSnl4yBOXd/nbX/8SVOcQJuxs9zk6uo2ls/GiNjMe2is5OZyhmefs3ZtcvvIwNJHNjSFVBsvMwPEpxc4VwrJi1CmYHH0IZatYo4NoMCqoKNF4ghFM2UOjAy1AHUWng8Gjqynzg/fYtyuK8XUecJF/fPrL4AIsJ2wOS86PP2x1RralhBmjWAFwnpPYJldh6xF+6clnWO7t8ZYEYt6hm19i8eGYbscimWduF4BBfB8TE5AoEbUVGA8awOaY2CGPgvMNhVR0zZJNmdA7f5/v//7z0DRgczg7Q0JFB4g0eMDS33rRaE0/NFhgc1+YznzyzKLh4F/+mQe++Dg2E5zC5Kdv88C1B5HCcjY7hTx1nSw6jDqCSCqrIonFvgGbkc1X7OQOJkdsUBNPP6A/P+TfvvV0yj+JMD3DhpqBdajWFMbgVRHMSCXO2cZTA4teOqdGh+C2oSmgtwEm8unnX+DqLz7OD29+yEerBcUjV6kWJ0iEoumgWlCZrC0rESRgehldH/DvXOexey5zdONNbHXMW//wN3D9NWgOoF5BgGFRUC8qOmLwGmmg9ST5i46AI2IzmEfSPwBSwrIG79OtzYTjH/07e/ffxyJ6ep/9LGcnY3AOiYY8pEMeb+1d7VPR8YdsbwzYPD2hGN/ijb/6Lif/+gp89A5kNSzO6OaCVhCbgAUiSgQy26FOs0+mQqAg4gGfp2pC04FgyUlrVjRQdsGMoL/H4Lt/wdR1k8cCdGtDRFhlefKkl7aIL9jxK46++jQsT0Cm4E9BVxBr8O0IwVqQpxYcEBRDAP4bbzlY8WiPuv8AAAAASUVORK5CYII="
             mask="url(#mask13100)"
             id="image13104" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,2993,10208)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13108"><tspan
             x="0 158.25027 204.85364"
             y="0"
             sodipodi:role="line"
             id="tspan13106">W:1</tspan></text>
        <g
           id="g13110">
          <path
             d="m 8739,6329 -85,-45 130,-40 z m -85,-45 130,-40 -85,-45 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13112" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46062,-0.8876,-0.8876,-0.46062,8655,6283)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#ff3f00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13116"><tspan
             x="0"
             y="0"
             id="tspan13114">E</tspan></text>
        <g
           id="g13118">
          <path
             d="m 3452,12558 v -479 l 2903,479 z m 0,-479 2903,479 v -479 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13120" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,3499,12376)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13124"><tspan
             x="0 111.81454 223.62909 270.23245 382.047 484.47382 531.07721 652.11182 782.53418 829.13757 922.3443 981.85577 1028.4591 1140.2737 1261.3083 1307.9116 1419.7262 1531.5408 1633.9675 1745.7821 1792.3855 1904.2001 2016.0146 2137.0493 2183.6526 2295.467 2407.2817 2565.532 2677.3464"
             y="0"
             sodipodi:role="line"
             id="tspan13122">EXISTING 4&quot; PRIVATE PVC SEWER</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,3502,12174)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13128"><tspan
             x="0 55.823456 158.25027 204.85364 316.66818 409.87491 530.90955 577.51294 689.32745 801.14203 922.17664 968.78003 1071.2068 1117.8102 1229.6248 1350.6594"
             y="0"
             sodipodi:role="line"
             id="tspan13126">(FIELD VERIFIED)</tspan></text>
        <g
           id="g13130">
          <path
             d="m 2457,11673 -107,-59 82,90 z"
             style="fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:#dd6e00;stroke-width:12.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13132" />
        </g>
        <path
           d="m 2444,11688 796,631 h 164"
           style="fill:none;stroke:#dd6e00;stroke-width:9;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13134" />
        <g
           id="g13136">
          <path
             d="m 5337,4744 -87,-46 203,-174 z m -87,-46 203,-174 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13138" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46402,-0.88582,-0.88582,-0.46402,5246,4708)"
           style="font-variant:normal;font-weight:normal;font-size:134.11px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00bfff;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13142"><tspan
             x="0 96.827736 134.11044"
             y="0"
             sodipodi:role="line"
             id="tspan13140">R/W</tspan></text>
        <g
           id="g13144">
          <path
             d="m 2685,16485 -89,-47 217,-197 z m -89,-47 217,-197 -89,-47 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13146" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46504,-0.88529,-0.88529,-0.46504,2595,16445)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13150"><tspan
             x="0 96.828171 186.28023"
             y="0"
             sodipodi:role="line"
             id="tspan13148">C&amp;G</tspan></text>
        <g
           id="g13152">
          <path
             d="m 6378,10323 v -278 l 861,278 z m 0,-278 861,278 v -278 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13154" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,6428,10141)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13158"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan13156">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,6741,10141)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13162"><tspan
             x="0 102.42682 223.46146 335.276"
             y="0"
             sodipodi:role="line"
             id="tspan13160">TREE</tspan></text>
        <g
           id="g13164">
          <path
             d="m 4999,9564 -116,-36 98,72 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13166" />
        </g>
        <path
           d="m 4990,9582 1177,602 h 163"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13168" />
        <g
           id="g13170">
          <path
             d="m 7981,7772 v -277 l 860,277 z m 0,-277 860,277 v -277 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13172" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,8031,7590)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13176"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan13174">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,8343,7590)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13180"><tspan
             x="0 102.42682 223.46146 335.276"
             y="0"
             sodipodi:role="line"
             id="tspan13178">TREE</tspan></text>
        <g
           id="g13182">
          <path
             d="m 6580,6560 -103,-64 77,94 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13184" />
        </g>
        <path
           d="m 6567,6575 1202,1058 h 164"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13186" />
        <g
           id="g13188">
          <path
             d="m 8656,5940 v -277 l 1613,277 z m 0,-277 1613,277 v -277 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13190" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,8705,5758)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13194"><tspan
             x="0 55.823456 167.638"
             y="0"
             sodipodi:role="line"
             id="tspan13192">(E)</tspan></text>
        <text
           xml:space="preserve"
           transform="matrix(1,0,0,-1,9020,5758)"
           style="font-variant:normal;font-weight:normal;font-size:167.638px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13198"><tspan
             x="0 158.25027 270.06482 372.49164 484.30618 605.34082 651.94415 763.75873 875.5733 996.60791 1089.8147"
             y="0"
             sodipodi:role="line"
             id="tspan13196">WATER VAULT</tspan></text>
        <g
           id="g13200">
          <path
             d="m 7782,6063 -102,66 118,-29 z"
             style="fill:#808080;fill-opacity:1;fill-rule:nonzero;stroke:#808080;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13202" />
        </g>
        <path
           d="m 7790,6081 654,-280 h 164"
           style="fill:none;stroke:#808080;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13204" />
        <g
           id="g13206">
          <path
             d="m 1138,14024 46,-88 39,133 z m 46,-88 39,133 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13208" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88296,0.46945,0.46945,-0.88296,1187,13940)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13212"><tspan
             x="0"
             y="0"
             id="tspan13210">S</tspan></text>
        <g
           id="g13214">
          <path
             d="m 6951,12734 46,-88 1687,998 z m 46,-88 1687,998 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13216" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.8852,0.46521,0.46521,-0.8852,7069,12685)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13220"><tspan
             x="0 89.452011 178.90402 216.18686 305.63889 387.58066 424.86353 521.69165 626.02997 663.31281 752.76483 842.2168 968.81757 1058.2695 1155.0977 1192.3805 1266.9462 1356.3982 1438.3401 1527.792 1624.6201 1714.0721"
             y="0"
             sodipodi:role="line"
             id="tspan13218">EXISTING SEWER LATERAL</tspan></text>
        <g
           id="g13222">
          <path
             d="m 8283,12376 46,-88 39,133 z m 46,-88 39,133 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13224" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88296,0.46945,0.46945,-0.88296,8332,12291)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13228"><tspan
             x="0"
             y="0"
             id="tspan13226">S</tspan></text>
        <g
           id="g13230">
          <path
             d="m 10834,13716 46,-87 39,132 z m 46,-87 39,132 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13232" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.8876,0.46062,0.46062,-0.8876,10883,13632)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13236"><tspan
             x="0"
             y="0"
             id="tspan13234">S</tspan></text>
        <g
           id="g13238">
          <path
             d="m 11744,15252 46,-88 39,132 z m 46,-88 39,132 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13240" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.8876,0.46062,0.46062,-0.8876,11792,15167)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13244"><tspan
             x="0"
             y="0"
             id="tspan13242">S</tspan></text>
        <g
           id="g13246">
          <path
             d="m 11187,14361 44,-85 65,142 z m 44,-85 65,142 44,-85 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13248" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88475,0.46606,0.46606,-0.88475,11230,14275)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13252"><tspan
             x="0"
             y="0"
             id="tspan13250">W</tspan></text>
        <g
           id="g13254">
          <path
             d="m 10733,16567 -88,-46 599,-927 z m -88,-46 599,-927 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13256" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.348525,-0.6641025,-0.88547,-0.4647,10668,16482)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13260"><tspan
             x="0 67.089134 134.17827 162.14046 229.2296 290.68607 318.64825 391.26947 469.52338 497.48557 553.40991 609.33429 645.04144 673.0036 740.09271 807.18188 879.8031 907.76526"
             y="0"
             sodipodi:role="line"
             id="tspan13258">EXISTING 16&quot; PVC W</tspan></text>
        <g
           id="g13262">
          <path
             d="m 9601,18600 -85,-45 143,-64 z m -85,-45 143,-64 -85,-45 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13264" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46606,-0.88475,-0.88475,-0.46606,9516,18557)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13268"><tspan
             x="0"
             y="0"
             id="tspan13266">W</tspan></text>
        <g
           id="g13270">
          <path
             d="m 4467,17073 -88,-46 133,-39 z m -88,-46 133,-39 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13272" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46945,-0.88296,-0.88296,-0.46945,4383,17024)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13276"><tspan
             x="0"
             y="0"
             id="tspan13274">S</tspan></text>
        <g
           id="g13278">
          <path
             d="m 5989,14175 -88,-46 531,-796 z m -88,-46 531,-796 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13280" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.3493575,-0.6636675,-0.88489,-0.46581,5910,14117)"
           style="font-variant:normal;font-weight:normal;font-size:134.112px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13284"><tspan
             x="0 67.08934 134.17868 162.14095 229.23029 290.68695 318.6492 391.27066 469.52478 497.48706 553.41162 589.11884 617.08112 684.17041 751.25977 823.88123 851.84351"
             y="0"
             sodipodi:role="line"
             id="tspan13282">EXISTING 8&quot; PVC S</tspan></text>
        <g
           id="g13286">
          <path
             d="m 10006,6528 -87,-46 132,-39 z m -87,-46 132,-39 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13288" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46062,-0.8876,-0.8876,-0.46062,9922,6479)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13292"><tspan
             x="0"
             y="0"
             id="tspan13290">S</tspan></text>
        <g
           id="g13294">
          <path
             d="m 3688,16593 -88,-46 515,-768 z m -88,-46 515,-768 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13296" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.348525,-0.6641025,-0.88547,-0.4647,3615,16524)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00dd00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13300"><tspan
             x="0 67.089134 134.17827 162.14046 229.2296 290.68607 318.64825 391.26947 469.52338 497.48557 553.40991 589.11707 617.07922 689.70044 756.78961 784.75177"
             y="0"
             sodipodi:role="line"
             id="tspan13298">EXISTING 3&quot; HP G</tspan></text>
        <g
           id="g13302">
          <path
             d="m 9071,6345 -88,-46 133,-39 z m -88,-46 133,-39 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13304" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46258,-0.88658,-0.88658,-0.46258,8983,6303)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00dd00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13308"><tspan
             x="0"
             y="0"
             id="tspan13306">G</tspan></text>
        <g
           id="g13310">
          <path
             d="m 5319,13487 -87,-46 132,-39 z m -87,-46 132,-39 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13312" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.47013,-0.8826,-0.8826,-0.47013,5231,13445)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00dd00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13316"><tspan
             x="0"
             y="0"
             id="tspan13314">G</tspan></text>
        <g
           id="g13318">
          <path
             d="m 4930,13579 -85,-45 130,-40 z m -85,-45 130,-40 -85,-44 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13320" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46945,-0.88296,-0.88296,-0.46945,4846,13533)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#ff3f00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13324"><tspan
             x="0"
             y="0"
             id="tspan13322">E</tspan></text>
        <g
           id="g13326">
          <path
             d="m 1816,16801 45,-85 65,143 z m 45,-85 65,143 44,-85 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13328" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88475,0.46606,0.46606,-0.88475,1860,16715)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13332"><tspan
             x="0"
             y="0"
             id="tspan13330">W</tspan></text>
        <g
           id="g13334">
          <path
             d="m 11282,8222 44,-85 65,142 z m 44,-85 65,142 45,-85 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13336" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88475,0.46606,0.46606,-0.88475,11325,8136)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13340"><tspan
             x="0"
             y="0"
             id="tspan13338">W</tspan></text>
        <g
           id="g13342">
          <path
             d="m 5433,5706 27,-92 91,127 z m 27,-92 91,127 27,-92 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13344" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.96123,0.27576,0.27576,-0.96123,5458,5614)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13348"><tspan
             x="0"
             y="0"
             id="tspan13346">W</tspan></text>
        <g
           id="g13350">
          <path
             d="m 10173,4848 46,-88 39,133 z m 46,-88 39,133 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13352" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88296,0.46945,0.46945,-0.88296,10222,4763)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13356"><tspan
             x="0"
             y="0"
             id="tspan13354">S</tspan></text>
        <g
           id="g13358">
          <path
             d="m 7623,3508 46,-88 39,133 z m 46,-88 39,133 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13360" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88296,0.46945,0.46945,-0.88296,7671,3423)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13364"><tspan
             x="0"
             y="0"
             id="tspan13362">S</tspan></text>
        <g
           id="g13366">
          <path
             d="m 6999,2447 46,-88 39,133 z m 46,-88 39,133 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13368" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88296,0.46945,0.46945,-0.88296,7048,2362)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13372"><tspan
             x="0"
             y="0"
             id="tspan13370">S</tspan></text>
        <path
           d="m 3708,8384 -14,26"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13374" />
        <path
           d="m 4239,8663 -14,26"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13376" />
        <path
           d="m 3821,8375 70,37"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13378" />
        <path
           d="m 4182,8565 -70,-37"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13380" />
        <g
           id="g13382">
          <path
             d="m 3814,8389 15,-28 -93,-30 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13384" />
        </g>
        <g
           id="g13386">
          <path
             d="m 4175,8579 15,-28 77,59 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13388" />
        </g>
        <g
           id="g13390">
          <path
             d="m 3927,8551 v -162 l 149,162 z m 0,-162 149,162 v -162 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13392" />
        </g>
        <path
           d="m 3997,8422 v 96 l -46,-64 h 69"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13394" />
        <path
           d="m 4052,8532 -5,-5 -4,5 4,4 5,-4 v -9 l -5,-9 -4,-5"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13396" />
        <path
           d="m 4748,9557 -57,109"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13398" />
        <path
           d="m 3938,9236 -14,27"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13400" />
        <path
           d="m 4648,9541 -188,-99"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13402" />
        <path
           d="m 4051,9228 188,99"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13404" />
        <g
           id="g13406">
          <path
             d="m 4641,9555 15,-28 77,59 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13408" />
        </g>
        <g
           id="g13410">
          <path
             d="m 4044,9242 15,-29 -93,-30 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13412" />
        </g>
        <g
           id="g13414">
          <path
             d="m 4275,9466 v -163 l 149,163 z m 0,-163 149,163 v -163 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13416" />
        </g>
        <path
           d="m 4354,9419 -4,9 -14,4 h -9 l -14,-4 -9,-14 -5,-23 v -23 l 5,-18 9,-9 14,-5 h 4 l 14,5 9,9 5,14 v 4 l -5,14 -9,9 -14,5 h -4 l -14,-5 -9,-9 -5,-14"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13418" />
        <path
           d="m 4400,9446 -5,-4 -4,4 4,5 5,-5 v -9 l -5,-9 -4,-5"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13420" />
        <path
           d="m 3711,9670 138,-263"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13422" />
        <path
           d="m 5680,10435 -56,107"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13424" />
        <path
           d="m 3892,9531 698,366"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13426" />
        <path
           d="m 5581,10418 -698,-366"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13428" />
        <g
           id="g13430">
          <path
             d="m 3884,9545 15,-28 -92,-31 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13432" />
        </g>
        <g
           id="g13434">
          <path
             d="m 5574,10432 14,-28 78,59 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13436" />
        </g>
        <g
           id="g13438">
          <path
             d="m 4626,10056 v -163 l 221,163 z m 0,-163 221,163 v -163 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13440" />
        </g>
        <path
           d="m 4650,10004 9,5 13,14 v -96"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13442" />
        <path
           d="m 4768,9927 v 96 l -45,-64 h 68"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13444" />
        <path
           d="m 4823,10036 -4,-4 -5,4 5,5 4,-5 v -9 l -4,-9 -5,-5"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13446" />
        <path
           d="m 4170,10426 34,-64"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13448" />
        <path
           d="m 3463,10142 -14,26"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13450" />
        <path
           d="m 4077,10397 -141,-74"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13452" />
        <path
           d="m 3576,10133 140,74"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13454" />
        <g
           id="g13456">
          <path
             d="m 4069,10411 15,-29 78,59 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13458" />
        </g>
        <g
           id="g13460">
          <path
             d="m 3568,10147 15,-28 -92,-30 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13462" />
        </g>
        <g
           id="g13464">
          <path
             d="m 3752,10346 v -162 l 148,162 z m 0,-162 148,162 v -162 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13466" />
        </g>
        <path
           d="m 3831,10313 h -46 l -4,-41 4,4 14,5 h 14 l 13,-5 9,-9 5,-14 v -9 l -5,-13 -9,-10 -13,-4 h -14 l -14,4 -4,5 -5,9"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13468" />
        <path
           d="m 3876,10327 -4,-5 -5,5 5,4 4,-4 v -10 l -4,-9 -5,-4"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13470" />
        <path
           d="m 2486,11355 -14,27"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13472" />
        <path
           d="m 2752,11495 -14,26"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13474" />
        <path
           d="m 2429,11258 -85,-45"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13476" />
        <path
           d="m 2865,11486 85,45 h 96"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13478" />
        <g
           id="g13480">
          <path
             d="m 2422,11272 15,-29 77,59 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13482" />
        </g>
        <g
           id="g13484">
          <path
             d="m 2857,11501 15,-29 -92,-30 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13486" />
        </g>
        <g
           id="g13488">
          <path
             d="m 3082,11612 v -162 l 148,162 z m 0,-162 148,162 v -162 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13490" />
        </g>
        <path
           d="m 3110,11556 v 5 l 5,9 4,4 10,5 h 18 l 9,-5 5,-4 4,-9 v -9 l -4,-10 -10,-13 -45,-46 h 64"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13492" />
        <path
           d="m 3206,11593 -4,-5 -5,5 5,4 4,-4 v -9 l -4,-10 -5,-4"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13494" />
        <path
           d="m 4213,7400 27,14"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13496" />
        <path
           d="m 4310,7215 27,14"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13498" />
        <path
           d="m 4115,7457 -44,85"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13500" />
        <path
           d="m 4302,7102 44,-85 h 96"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13502" />
        <g
           id="g13504">
          <path
             d="m 4130,7464 -29,-15 59,-77 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13506" />
        </g>
        <g
           id="g13508">
          <path
             d="m 4316,7110 -29,-15 -30,92 z"
             style="fill:#ff0000;fill-opacity:1;fill-rule:nonzero;stroke:#ff0000;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13510" />
        </g>
        <g
           id="g13512">
          <path
             d="m 4478,7098 v -162 l 131,162 z m 0,-162 131,162 v -162 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13514" />
        </g>
        <path
           d="m 4502,7047 9,5 14,13 v -96"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13516" />
        <path
           d="m 4585,7079 -5,-5 -5,5 5,5 5,-5 v -9 l -5,-9 -5,-5"
           style="fill:none;stroke:#ff0000;stroke-width:12;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
           id="path13518" />
        <g
           id="g13520">
          <path
             d="m 8552,16072 -112,-59 693,-1049 z m -112,-59 693,-1049 -111,-58 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13522" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.3486525,-0.664035,-0.88538,-0.46487,8494,15973)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13526"><tspan
             x="0 67.089088 134.17818 162.14035 229.22945 290.68585 318.64804 391.2692 469.52304 497.48523 553.40955 589.11664 617.0788 684.16791 712.13007 745.62433 812.71344 879.80249 946.8916 1019.5128 1092.1339"
             y="0"
             sodipodi:role="line"
             id="tspan13524">EXISTING 6&quot; S (ABAND)</tspan></text>
        <g
           id="g13528">
          <path
             d="m 9079,16822 -88,-46 686,-1093 z m -88,-46 686,-1093 -88,-46 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13530" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.46504,-0.88529,-0.88529,-0.46504,8996,16771)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#0000ff;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13534"><tspan
             x="0 74.565735 149.13147 174.74669 212.02956 308.85773 398.30978 435.59265 525.04474 614.49677 711.32495 748.60785 860.32233 949.77435 1046.6025 1083.8854 1173.3375"
             y="0"
             sodipodi:role="line"
             id="tspan13532">10' RAISED MEDIAN</tspan></text>
        <g
           id="g13536">
          <path
             d="m 9308,12915 46,-88 1687,998 z m 46,-88 1687,998 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13538" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.8852,0.46521,0.46521,-0.8852,9426,12866)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13542"><tspan
             x="0 89.452011 178.90402 216.18686 305.63889 387.58066 424.86353 521.69165 626.02997 663.31281 752.76483 842.2168 968.81757 1058.2695 1155.0977 1192.3805 1266.9462 1356.3982 1438.3401 1527.792 1624.6201 1714.0721"
             y="0"
             sodipodi:role="line"
             id="tspan13540">EXISTING SEWER LATERAL</tspan></text>
        <g
           id="g13544">
          <path
             d="m 2838,14917 46,-88 1687,999 z m 46,-88 1687,999 47,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13546" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.8852,0.46521,0.46521,-0.8852,2956,14869)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13550"><tspan
             x="0 89.452011 178.90402 216.18686 305.63889 387.58066 424.86353 521.69165 626.02997 663.31281 752.76483 842.2168 968.81757 1058.2695 1155.0977 1192.3805 1266.9462 1356.3982 1438.3401 1527.792 1624.6201 1714.0721"
             y="0"
             sodipodi:role="line"
             id="tspan13548">EXISTING SEWER LATERAL</tspan></text>
        <g
           id="g13552">
          <path
             d="m 3461,17667 46,-88 1687,999 z m 46,-88 1687,999 47,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13554" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88538,0.46487,0.46487,-0.88538,3582,17620)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13558"><tspan
             x="0 89.452118 178.90424 216.18713 305.63925 387.58115 424.86404 521.69226 626.0307 663.3136 789.91455 879.36664 961.30853 1050.7606 1147.5889 1184.8718 1259.4376 1348.8896 1430.8315 1520.2837 1617.1119 1706.5641"
             y="0"
             sodipodi:role="line"
             id="tspan13556">EXISTING WATER LATERAL</tspan></text>
        <g
           id="g13560">
          <path
             d="m 8790,6906 46,-88 1688,999 z m 46,-88 1688,999 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13562" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88515,0.4653,0.4653,-0.88515,8911,6859)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#00a5dd;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13566"><tspan
             x="0 89.451797 178.90359 216.18636 305.63815 387.57974 424.86252 521.69037 626.02844 663.31122 789.91168 879.36346 961.30505 1050.7568 1147.5847 1184.8676 1259.433 1348.8848 1430.8264 1520.2782 1617.1061 1706.5579"
             y="0"
             sodipodi:role="line"
             id="tspan13564">EXISTING WATER LATERAL</tspan></text>
        <g
           id="g13568">
          <path
             d="m 8769,4111 47,-88 1687,998 z m 47,-88 1687,998 46,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13570" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.8852,0.46521,0.46521,-0.8852,8887,4062)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13574"><tspan
             x="0 89.452011 178.90402 216.18686 305.63889 387.58066 424.86353 521.69165 626.02997 663.31281 752.76483 842.2168 968.81757 1058.2695 1155.0977 1192.3805 1266.9462 1356.3982 1438.3401 1527.792 1624.6201 1714.0721"
             y="0"
             sodipodi:role="line"
             id="tspan13572">EXISTING SEWER LATERAL</tspan></text>
        <g
           id="g13576">
          <path
             d="m 10433,4251 47,-87 38,132 z m 47,-87 38,132 47,-88 z"
             style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:12.5;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-opacity:1"
             id="path13578" />
        </g>
        <text
           xml:space="preserve"
           transform="matrix(0.88992,0.45611,0.45611,-0.88992,10482,4167)"
           style="font-variant:normal;font-weight:normal;font-size:134.111px;font-family:Arial;-inkscape-font-specification:ArialMT;writing-mode:lr-tb;fill:#dd6e00;fill-opacity:1;fill-rule:nonzero;stroke:none"
           id="text13582"><tspan
             x="0"
             y="0"
             id="tspan13580">S</tspan></text>
      </g>
    </g>
  </g>
</svg>
